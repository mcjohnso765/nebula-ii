* NGSPICE file created from team_07_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

.subckt team_07_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[3] la_oenb[4]
+ la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
X_05903_ _01585_ net122 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__nand2_2
X_10932__582 vssd1 vssd1 vccd1 vccd1 _10932__582/HI net582 sky130_fd_sc_hd__conb_1
X_09671_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\] _04725_ net1170
+ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a21oi_1
X_06883_ net108 _02550_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__nor2_1
XANTENNA__07534__B2 _02119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ net457 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__nand2b_1
X_05834_ _01505_ _01511_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08553_ net139 _04005_ _03963_ vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__o21ai_1
X_05765_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\]
+ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout162_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07504_ _00759_ _01610_ net100 vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__a21o_1
X_08484_ _03817_ _03898_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_18_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05696_ _01318_ _01393_ _01394_ _01408_ vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__a31o_2
XFILLER_0_43_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07435_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] _03014_
+ net479 vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07366_ net967 _02965_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09105_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ _04342_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__a21o_1
X_06317_ _01970_ _01971_ _01972_ _01992_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__and4_1
XFILLER_0_116_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07065__A3 _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07297_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09036_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ _04291_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06248_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] net183 vssd1 vssd1
+ vccd1 vccd1 _01925_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold340 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06179_ net279 net159 net147 net281 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__o22a_1
Xhold351 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_right vssd1
+ vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold373 team_07_WB.instance_to_wrap.team_07.label_num_bus\[2\] vssd1 vssd1 vccd1
+ vccd1 net1043 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold384 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[3\] vssd1 vssd1
+ vccd1 vccd1 net1054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[5\] vssd1
+ vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06576__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ net465 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
XANTENNA__06411__B _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09869_ _04866_ _04867_ net1091 net241 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_29_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07856__A1_N _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10829__505 vssd1 vssd1 vccd1 vccd1 _10829__505/HI net505 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_103_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07828__A2 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10713_ clknet_leaf_60_wb_clk_i _00544_ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10644_ clknet_leaf_41_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[1\]
+ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10575_ clknet_leaf_24_wb_clk_i _00443_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07461__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06602__A net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08961__A0 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output56_A net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07516__A1 _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10009_ clknet_leaf_33_wb_clk_i _00006_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05550_ _01259_ _01261_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08963__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05481_ _00965_ _01175_ _01193_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__and3_2
XFILLER_0_11_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07220_ _02864_ _02866_ _02869_ _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__o31a_1
XFILLER_0_129_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07151_ net168 _02033_ _02775_ _02803_ _02773_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a32o_1
XFILLER_0_125_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10091__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06055__Y _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06102_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\]
+ _01784_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__nor3_1
XANTENNA__06255__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05400__B _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07082_ _01618_ net253 _02735_ _02127_ _02734_ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a221o_2
XANTENNA__06255__B2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06033_ net197 net185 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__nand2_2
XFILLER_0_112_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout105 _01691_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_4
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06558__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout116 net117 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__buf_2
XANTENNA__08952__B1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout127 net128 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout138 _01648_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_4
Xfanout149 net150 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_4
X_07984_ _01700_ _01732_ _03375_ _03526_ _03405_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__a41o_1
X_09723_ net250 _04761_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_52_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06935_ _02501_ _02591_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__nor2_1
XANTENNA__07507__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_87_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07507__B2 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09654_ _04711_ _04712_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__nor2_2
X_06866_ net286 net434 _02483_ _02536_ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08605_ _01242_ _01248_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05817_ _01496_ _01510_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__nor2_1
X_09585_ _04667_ _04668_ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__nor2_1
X_06797_ _00696_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1
+ vccd1 vccd1 _02468_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout165_X net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07062__B _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08536_ _03976_ _03990_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05748_ net1108 _01445_ _01447_ _00787_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[8\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10179__RESET_B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05679_ _01347_ _01350_ _01366_ _01391_ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__o211a_1
X_08467_ net460 _03936_ _03937_ _03938_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__o32a_1
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07418_ _03004_ _03005_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[12\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08398_ _03709_ _03872_ _03850_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__o21a_1
XANTENNA__05150__X _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07349_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[14\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[13\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[12\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[15\] vssd1 vssd1
+ vccd1 vccd1 _02958_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05310__B _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10360_ clknet_leaf_22_wb_clk_i net727 net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.rand_num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09019_ net251 _04279_ _04281_ net403 net876 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__a32o_1
X_10291_ clknet_leaf_45_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[4\]
+ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold170 _00498_ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06422__A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold181 team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[0\] vssd1 vssd1 vccd1
+ vccd1 net851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06549__A2 _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07237__B _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06721__A2 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08067__A_N net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06485__A1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06485__B2 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10627_ clknet_leaf_49_wb_clk_i _00491_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05220__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10558_ clknet_leaf_19_wb_clk_i _00426_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06603__Y _02276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489_ clknet_leaf_14_wb_clk_i _00357_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08023__S _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06051__B net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04981_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
X_06720_ _01675_ _02021_ net258 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06651_ _02321_ _02322_ _02323_ _02178_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a31o_1
X_05602_ net443 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\] vssd1 vssd1
+ vccd1 vccd1 _01315_ sky130_fd_sc_hd__nand2_2
X_09370_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ _04530_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__a31o_1
X_06582_ _02196_ _02245_ _02246_ net84 _02255_ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05533_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right net424
+ net423 _01206_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__o221a_1
X_08321_ _03715_ _03798_ _03752_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08252_ _01281_ _01303_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__nand2_1
X_05464_ _00966_ _01103_ _01107_ _01112_ _01176_ vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07203_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[7\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\]
+ net449 vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08183_ _03655_ _03660_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__or2_2
XFILLER_0_43_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09414__A1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05395_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ _00795_ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__or2_2
XFILLER_0_131_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07134_ _02785_ _02786_ _02787_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07065_ _01679_ _01904_ _01936_ _02687_ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__o41a_1
XFILLER_0_113_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06016_ net181 net172 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__or2_4
XFILLER_0_100_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05451__A2 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07189__C1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06400__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ _03415_ _03521_ _03486_ _03519_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__or4b_1
XFILLER_0_57_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09706_ _04750_ _04751_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\]
+ _04730_ vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__a2bb2o_1
X_06918_ _02512_ _02516_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__nor2_1
XANTENNA__08169__A net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ _03374_ _03382_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__nor2_1
X_09637_ net958 _04700_ _04701_ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__a21o_1
X_06849_ net262 _02509_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__nor2_1
X_09568_ net480 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ _04657_ _04658_ vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08519_ _03981_ _03982_ vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__nor2_1
XANTENNA__10755__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09499_ _00667_ _04626_ net290 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06467__A1 _02060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07520__B _02744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06219__A1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ clknet_leaf_23_wb_clk_i _00303_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05975__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10343_ clknet_leaf_56_wb_clk_i _00283_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05978__B1 _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10274_ clknet_leaf_73_wb_clk_i _00266_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout480 net484 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout491 net492 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09341__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06046__B _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05180_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00890_ vssd1 vssd1
+ vccd1 vccd1 _00893_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09966__RESET_B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07610__A1_N _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08870_ net445 net808 net246 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08383__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07821_ _03371_ _03375_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__nor2_1
X_04964_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\] vssd1
+ vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
X_07752_ _03303_ _03306_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__nand2_1
X_06703_ _02066_ _02362_ net83 _02079_ _02236_ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__a221o_1
XANTENNA__10453__RESET_B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ _01678_ _01903_ _01935_ _03174_ _01905_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__a311o_1
X_09422_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\] _04567_
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[2\] vssd1
+ vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a31o_1
XANTENNA__07894__A0 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06697__B2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06634_ _02304_ _02306_ _02178_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a21o_1
X_09353_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ _04520_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06565_ _02218_ _02225_ _02233_ _02238_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout242_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08304_ _03702_ _03778_ _03779_ _03780_ _03711_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__a41o_1
X_05516_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ _01223_ _01228_ _01199_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__a211o_1
X_09284_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06496_ _01620_ net274 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__nor2_2
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08235_ _03674_ _03712_ _03713_ net477 vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__o211a_1
X_05447_ _01060_ _01089_ _01048_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout128_X net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08166_ _00704_ _03647_ _00703_ vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_95_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05378_ _00969_ _01083_ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__nor2_2
XANTENNA__07949__B2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07117_ net95 _02770_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08097_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[13\]
+ _00814_ net483 vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06082__C1 _01748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07048_ _02363_ _02366_ _02702_ _02697_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__o31a_1
XANTENNA__06621__A1 _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input2_X net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _04258_ _04260_ _04267_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10961_ net602 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XANTENNA__06137__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10892_ net649 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_39_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06147__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05986__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06434__X _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__B2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06612__A1 _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10326_ clknet_leaf_51_wb_clk_i _00044_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ clknet_leaf_75_wb_clk_i _00249_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10188_ clknet_leaf_82_wb_clk_i net712 net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06679__A1 _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06609__X _02282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06350_ _00710_ net215 net177 _01723_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08971__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05301_ net431 _00999_ vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_20_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06281_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] net133 _01934_ _01938_
+ net262 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_115_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05232_ _00899_ net300 _00944_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08020_ net866 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__nand2_1
XANTENNA__05896__A _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08272__A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05163_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00876_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08053__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06504__B _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05094_ _00809_ _00818_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__or2_1
X_09971_ clknet_leaf_83_wb_clk_i _00076_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08922_ net241 _04230_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09553__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ net455 net413 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ _04187_ vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__o31a_1
XFILLER_0_23_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06520__A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06906__A2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07804_ _03351_ _03350_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__nand2b_1
X_08784_ _04139_ _04140_ net195 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__a21oi_1
X_05996_ net134 net123 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__nand2_8
XANTENNA__05136__A team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07735_ net285 _01105_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04947_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\] vssd1
+ vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07666_ net126 net141 _02260_ _02768_ _01729_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__a32o_1
XFILLER_0_48_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07331__A2 _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ net481 _04561_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06617_ _01625_ _02140_ _02289_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07597_ _03152_ _03154_ _03155_ _03151_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__o31a_1
XFILLER_0_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout245_X net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10862__538 vssd1 vssd1 vccd1 vccd1 _10862__538/HI net538 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_138_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09336_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__nand3_1
XFILLER_0_118_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06548_ net287 _00748_ _02180_ net85 net266 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07501__D _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07095__A1 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09267_ net336 _04426_ _04464_ net900 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06479_ _02034_ _02035_ _02038_ _02152_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a31o_2
XFILLER_0_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06842__A1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08218_ net459 _03693_ _03696_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ _04369_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__nand3_1
XFILLER_0_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08149_ net475 _03634_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_112_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08910__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10111_ clknet_leaf_36_wb_clk_i _00149_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08347__A1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10042_ _00062_ _00640_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__07526__A _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09544__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold63 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[5\] vssd1
+ vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 _00115_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10944_ team_07_WB.instance_to_wrap.audio vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_27_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10323__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06530__B1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10875_ net551 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XFILLER_0_112_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05884__A2 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_85_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07086__A1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06605__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_5 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10309_ clknet_leaf_45_wb_clk_i net804 net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05850_ _01534_ _01537_ _01540_ _01541_ _01536_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__a41o_1
XANTENNA__08966__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05781_ _01461_ _01462_ _01463_ _01464_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__and4b_1
X_07520_ _01873_ _02744_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__or2_2
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07451_ net453 net413 vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__and2_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06521__B1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06402_ _02060_ _02071_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__nand2_1
X_07382_ net1163 _02981_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09121_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ _04355_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06333_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _01631_ _02007_
+ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_40_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06285__C1 _01961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06264_ net180 _01923_ _01925_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09052_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ _04304_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06074__X _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05215_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ _00897_ _00915_ _00927_ vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__a311o_1
X_08003_ _03552_ _03553_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__xnor2_1
Xhold500 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[8\] vssd1 vssd1
+ vccd1 vccd1 net1170 sky130_fd_sc_hd__dlygate4sd3_1
X_06195_ _01855_ _01872_ _01875_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__o21ai_1
Xhold511 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05146_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[5\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[7\]
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] vssd1 vssd1 vccd1 vccd1
+ _00859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10815__RESET_B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09954_ clknet_leaf_90_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[3\]
+ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_38_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05077_ net426 _00694_ net434 _00675_ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08905_ _01405_ net441 net440 vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__or3b_1
X_09885_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\] _01773_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__o21ai_1
X_08836_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\] _04142_
+ net875 vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07552__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10346__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08767_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] net805 net235 vssd1
+ vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__mux2_1
X_05979_ _01647_ _01655_ _01672_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07718_ _01590_ _01598_ _01065_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08698_ _00693_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ _01238_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_64_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07081__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07649_ _03204_ _03206_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10660_ clknet_leaf_3_wb_clk_i _00515_ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_82_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06128__C net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09319_ _00661_ _04500_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10591_ clknet_leaf_38_wb_clk_i _00455_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XANTENNA__07240__A1 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05983__B net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06043__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
XANTENNA__07240__B2 _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput75 net391 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_0_37_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10025_ clknet_leaf_53_wb_clk_i _00002_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10927_ net577 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10884__560 vssd1 vssd1 vccd1 vccd1 _10884__560/HI net560 sky130_fd_sc_hd__conb_1
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05223__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10858_ net534 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_39_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10789_ clknet_leaf_76_wb_clk_i _00610_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06806__A1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05000_ net12 net11 net14 net13 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__or4_1
XANTENNA__06054__B net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10297__RESET_B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09508__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07782__A2 _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06951_ _02506_ _02508_ net174 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05902_ _01585_ net121 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _01763_ _04712_ _04721_ _04726_ vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__a31o_1
X_06882_ net116 _02478_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08621_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__nand2_1
X_05833_ _01506_ _01520_ _01523_ _01525_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_85_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08552_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[7\]
+ _03611_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__xor2_1
X_05764_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\]
+ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_89_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07503_ _03058_ _03061_ _03062_ _03050_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.stageDetect
+ sky130_fd_sc_hd__o31a_1
XANTENNA__05414__A team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ net468 net474 _03640_ _03659_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_18_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05695_ net491 _01404_ _01407_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__or3_1
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07434_ _03014_ _03015_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[18\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07365_ _02965_ _02972_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_sck_rs_enable
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout322_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09104_ net212 _04344_ _04345_ net399 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06316_ _01983_ _01991_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06245__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07296_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09035_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ _04291_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout110_X net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06247_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] net173 _01923_ vssd1
+ vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold330 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] vssd1 vssd1
+ vccd1 vccd1 net1000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[1\] vssd1
+ vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__dlygate4sd3_1
X_06178_ net281 net147 _01858_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__a21oi_1
Xhold352 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_right vssd1
+ vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold363 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold374 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_select
+ vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__dlygate4sd3_1
X_05129_ _00837_ _00838_ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold385 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\] vssd1 vssd1
+ vccd1 vccd1 net1055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07076__A _02726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09937_ net466 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
XANTENNA__06411__C net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09868_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ _04228_ net263 vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_29_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911__656 vssd1 vssd1 vccd1 vccd1 net656 _10911__656/LO sky130_fd_sc_hd__conb_1
X_08819_ _04166_ _04167_ _04144_ vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09799_ net1023 _04808_ _04819_ vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__a21o_1
X_10868__544 vssd1 vssd1 vccd1 vccd1 _10868__544/HI net544 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_103_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ clknet_leaf_71_wb_clk_i _00543_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10643_ clknet_leaf_41_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[0\]
+ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10574_ clknet_leaf_24_wb_clk_i _00442_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09450__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05472__B1 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10390__RESET_B net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06602__B _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07516__A2 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07714__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ clknet_leaf_55_wb_clk_i _00005_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07348__A1_N net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05480_ _00964_ _01109_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07150_ net150 net129 _01710_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06101_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[19\] _01783_
+ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__or2_2
X_07081_ net95 net93 net88 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06032_ net200 net189 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__nor2_4
XANTENNA__06352__X _02027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout106 _01651_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout117 _01608_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_4
Xfanout128 _01594_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_4
Xfanout139 net140 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
X_07983_ _00746_ _03354_ _03363_ net267 vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__o22a_1
X_09722_ _04731_ _04760_ _04762_ _04730_ net998 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__a32o_1
XANTENNA__05128__B team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06934_ net433 _01652_ _01700_ _02503_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_52_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07507__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ net1029 _04711_ _04713_ _04715_ vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__a22o_1
X_06865_ net282 _02474_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_2_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout272_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08604_ _01243_ _01758_ _04035_ _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__nand4_2
X_05816_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] _01486_
+ _01490_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__a21oi_1
X_09584_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\] _04665_ net1058
+ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06191__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06796_ _00695_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1
+ vccd1 vccd1 _02467_ sky130_fd_sc_hd__nor2_2
XFILLER_0_132_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06191__B2 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05144__A team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08535_ _03974_ _03990_ _03978_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__a21o_1
X_05747_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\]
+ _01446_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__and3_1
XANTENNA__07062__C _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10980__621 vssd1 vssd1 vccd1 vccd1 _10980__621/HI net621 sky130_fd_sc_hd__conb_1
XFILLER_0_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout158_X net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08466_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] net460
+ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__nand2_1
X_05678_ _01345_ _01378_ _01390_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07417_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\] _03003_
+ net233 vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07691__B2 _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03804_ _03847_
+ _00727_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__o31a_1
XFILLER_0_80_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ net490 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _02956_
+ _02957_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing_mod_locator.nxt_mod_row
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_122_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10148__RESET_B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07279_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09018_ _04280_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10290_ clknet_leaf_45_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[3\]
+ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold160 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[6\] vssd1 vssd1
+ vccd1 vccd1 net841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[14\] vssd1 vssd1
+ vccd1 vccd1 net852 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06422__B net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[21\]
+ vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06706__B1 _02235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05989__A _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07540__Y _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07682__A1 _02699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10626_ clknet_leaf_49_wb_clk_i net897 net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05995__Y _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10557_ clknet_leaf_19_wb_clk_i _00425_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05445__B1 _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10488_ clknet_leaf_25_wb_clk_i _00356_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07198__B1 _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04980_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06650_ _02107_ _02295_ _02308_ _02139_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a22oi_1
XANTENNA__08974__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10964__605 vssd1 vssd1 vccd1 vccd1 _10964__605/HI net605 sky130_fd_sc_hd__conb_1
XFILLER_0_87_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05601_ _01300_ _01313_ _01280_ _01297_ vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__o211a_1
X_06581_ _02231_ _02253_ _02254_ _02248_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08320_ net465 _03784_ _03796_ _03797_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__o22a_1
X_05532_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ _01231_ _01244_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07122__B1 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__RESET_B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08251_ _03685_ _03727_ _03728_ _01384_ net461 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07673__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05463_ _01100_ _01105_ _01111_ _01048_ vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_31_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07202_ _02827_ _02844_ _02847_ net167 _02853_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[2\]
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08182_ net474 net473 vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05394_ _01000_ net191 _01019_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__or3_2
XFILLER_0_42_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07133_ _02754_ _02773_ _02781_ _02733_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout118_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07178__X _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07064_ net129 _01904_ _01936_ _02684_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06523__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06015_ net181 net172 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07189__B1 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout487_A team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06400__A2 _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07966_ net281 net109 net275 _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__o31a_1
X_09705_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\] _04749_ _04731_
+ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06917_ _02579_ _02586_ _02587_ _02578_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a31o_1
X_07897_ _03451_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09636_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[20\] _04698_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__and3b_1
X_06848_ _02518_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09567_ _04657_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ _04548_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_136_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06779_ net182 _02447_ _02449_ _02450_ _02432_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08518_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\]
+ _03979_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07801__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09498_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] vssd1
+ vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08449_ _03632_ _03662_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nand2_1
XANTENNA__07664__A1 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07664__B2 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08861__B1 _01748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05321__B _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10411_ clknet_leaf_23_wb_clk_i _00302_ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_104_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05427__B1 _01104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10342_ clknet_leaf_54_wb_clk_i _00282_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_115_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05978__A1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06433__A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10273_ clknet_leaf_73_wb_clk_i _00265_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout90_X net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10917__662 vssd1 vssd1 vccd1 vccd1 net662 _10917__662/LO sky130_fd_sc_hd__conb_1
XFILLER_0_100_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_39_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout470 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[2\] vssd1
+ vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_2
Xfanout481 net483 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_2
Xfanout492 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_2
XFILLER_0_45_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08852__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10609_ clknet_leaf_47_wb_clk_i _00473_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08969__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06062__B team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07820_ _03372_ _03374_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__nor2_1
X_07751_ _03304_ _03305_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__or2_1
X_04963_ net53 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
XANTENNA__09332__A1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06702_ net115 net111 _02148_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07682_ _02699_ _03238_ _03239_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_126_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09421_ _04571_ _04573_ _04574_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__and3_1
X_06633_ _02119_ _02289_ _02305_ _02165_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__o22a_1
XANTENNA__07902__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ _04520_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__a21oi_1
X_06564_ _02160_ net85 _02214_ _02237_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a31o_1
XANTENNA__06518__A _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08303_ _03702_ _03778_ _03779_ _03780_ _03711_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a41oi_1
XFILLER_0_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05515_ net424 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__nor2_1
X_09283_ _04475_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__inv_2
X_06495_ _02119_ _02168_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout235_A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08234_ _00711_ team_07_WB.instance_to_wrap.team_07.lcdOutput.modSquaresPixel team_07_WB.instance_to_wrap.team_07.lcdOutput.modHighlightPixel
+ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__or3b_2
X_05446_ _01086_ _01096_ _01078_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08165_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\] _03647_
+ vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout402_A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05377_ _00966_ _01050_ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07116_ net278 net86 net93 vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08096_ _03600_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[13\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06082__B1 _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload80 clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__inv_12
X_07047_ _02065_ net84 _02692_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__and3_1
XANTENNA__06621__A2 _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04264_ _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__nor4_1
XANTENNA__07582__B1 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ _01692_ _03319_ _03491_ _03492_ net106 vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__o32a_1
XFILLER_0_138_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10960_ net601 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_98_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07334__A0 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\] _04688_ vssd1
+ vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__or2_1
XANTENNA__06688__A2 _01413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07885__A1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ net648 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_70_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10011__Q team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07090__Y _02744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07637__A1 _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07637__B2 _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10163__RESET_B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05986__B net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10325_ clknet_leaf_54_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[2\]
+ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06612__A2 _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ clknet_leaf_75_wb_clk_i _00248_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_10187_ clknet_leaf_82_wb_clk_i net697 net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07722__A _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06679__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06338__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07628__A1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05300_ _00996_ _01005_ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06280_ _01933_ _01947_ _01953_ _01956_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05231_ net449 _00840_ net398 _00832_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05162_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00875_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05093_ _00809_ _00818_ vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__nor2_1
X_09970_ clknet_leaf_82_wb_clk_i _00075_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[19\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05406__A3 _01104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08921_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[2\]
+ _04228_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08852_ net451 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ net297 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ _04186_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07803_ _01102_ net112 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__or2_1
X_08783_ _01454_ _04143_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05995_ net132 net127 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout185_A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07734_ net279 _01104_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__nor2_1
X_04946_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1 vssd1 vccd1
+ vccd1 _00686_ sky130_fd_sc_hd__inv_2
XANTENNA__06119__A1 _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10674__RESET_B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07665_ _01811_ _02055_ _03081_ _03222_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout352_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[7\]
+ _04560_ _04559_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06616_ _02265_ _02288_ _02272_ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07596_ _02082_ _03079_ _03100_ _02744_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_66_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06248__A team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09335_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_138_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06547_ net266 net84 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_138_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout140_X net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09266_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ net336 _04459_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__and4_1
XFILLER_0_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06478_ net187 net181 _02151_ _01684_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_62_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06535__X _02209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08217_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel _01296_
+ _03694_ _03695_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__a2bb2o_1
X_10903__569 vssd1 vssd1 vccd1 vccd1 _10903__569/HI net569 sky130_fd_sc_hd__conb_1
X_05429_ _01020_ _01053_ _01068_ vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__a21oi_1
X_09197_ net404 _04375_ _04412_ vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ net475 _03634_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08079_ _03592_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10110_ clknet_leaf_60_wb_clk_i team_07_WB.instance_to_wrap.team_07.boomGen.boomDetect
+ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.boomGen.boomPixel
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout98_A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10041_ _00061_ _00639_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__07526__B net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 _00112_ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[23\]
+ vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10943_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_cs vssd1 vssd1
+ vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10874_ net550 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XANTENNA__05333__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05997__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07086__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06445__X _02119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06605__B _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08035__A1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08035__B2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_54_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10308_ clknet_leaf_44_wb_clk_i net745 net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_10239_ clknet_leaf_82_wb_clk_i net690 net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05780_ _01465_ _01478_ net478 _01422_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10085__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07849__B2 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07450_ net455 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06521__B2 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06401_ _02074_ _02060_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_44_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07381_ _02974_ _02981_ _02982_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[5\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09120_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ _04355_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__or2_1
X_06332_ net289 _00754_ net87 net101 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09051_ net251 _04303_ _04304_ net407 net1136 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_13_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06263_ _01649_ _01938_ _01939_ _01934_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08002_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__xor2_1
X_05214_ _00918_ _00926_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08026__A1 _00706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold501 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06194_ _01716_ net102 _01873_ _01874_ _01683_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__o311a_1
XFILLER_0_12_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06037__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold512 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[2\] vssd1 vssd1
+ vccd1 vccd1 net1182 sky130_fd_sc_hd__dlygate4sd3_1
X_05145_ _00855_ _00856_ _00857_ vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout100_A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07186__X _02838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09953_ clknet_leaf_84_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[2\]
+ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_05076_ net431 _00695_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] _00674_
+ _00799_ vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_38_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08904_ net1053 _04217_ net264 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__o21a_1
X_09884_ net1092 net153 net151 _04877_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__a22o_1
X_08835_ _04176_ _04177_ net196 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout188_X net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] net820 net234 vssd1
+ vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__mux2_1
X_05978_ net163 _01669_ _01664_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07717_ _01649_ _01667_ _01743_ _03270_ _03272_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.borderGen.synchronized_rectangle_pixel
+ sky130_fd_sc_hd__a41o_1
X_04929_ net435 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
X_08697_ _00693_ _01238_ _01242_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07081__B net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07648_ net135 net128 _01743_ _03205_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_64_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07579_ _03130_ _03133_ _03134_ _03137_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__or4_1
XFILLER_0_75_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09318_ _00661_ net333 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08265__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ clknet_leaf_38_wb_clk_i _00454_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09249_ net230 _04451_ _04452_ net406 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07537__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XANTENNA__06441__A _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05787__C1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10024_ clknet_leaf_42_wb_clk_i net1009 net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input30_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10440__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10926_ net576 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05998__Y _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10857_ net533 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_2_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10788_ clknet_leaf_12_wb_clk_i _00609_ net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06019__B1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08042__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06351__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06950_ net433 net145 _02620_ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a21o_1
XANTENNA__08977__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05901_ _01579_ _01581_ _01584_ _01587_ _01593_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__a41o_1
XFILLER_0_94_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06881_ net116 _02478_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08620_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04046_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__and3_1
X_05832_ _01506_ _01520_ _01523_ _01525_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08551_ net146 _03652_ _03996_ _04004_ vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_85_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05763_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\]
+ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__nor4b_1
X_07502_ _02352_ _03060_ _03059_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08482_ net467 _03637_ _03641_ _03819_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__o31ai_1
X_05694_ _01402_ _01406_ net438 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07433_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\] _03013_
+ net233 vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout148_A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07364_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\] _02970_
+ _02971_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__or3b_1
XFILLER_0_116_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09444__B1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09103_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ _04342_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06315_ _01974_ _01984_ _01990_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07295_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09034_ net252 _04290_ _04292_ net405 net1067 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__a32o_1
X_06246_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] net183 vssd1 vssd1
+ vccd1 vccd1 _01923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold320 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[17\]
+ vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06177_ net285 net161 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__nor2_1
Xhold331 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_up vssd1
+ vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout103_X net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 _00027_ vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\] vssd1 vssd1 vccd1
+ vccd1 net1023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_left vssd1
+ vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__dlygate4sd3_1
X_05128_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__nand2_1
Xhold375 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10313__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold386 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05059_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\] _00788_ vssd1
+ vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__or2_1
X_09936_ net466 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09867_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ _04228_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_107_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06725__A1_N _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\] _01448_
+ _04160_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__or3_1
XANTENNA__06194__C1 _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09798_ _04818_ _04811_ _04817_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__and3b_1
XANTENNA__07930__B1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08749_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ net238 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10711_ clknet_leaf_68_wb_clk_i _00542_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06497__B1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10909__575 vssd1 vssd1 vccd1 vccd1 _10909__575/HI net575 sky130_fd_sc_hd__conb_1
XFILLER_0_36_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10642_ clknet_leaf_45_wb_clk_i net888 net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06436__A _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10573_ clknet_leaf_25_wb_clk_i _00441_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07461__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06171__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06421__B1 _02080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10007_ clknet_leaf_42_wb_clk_i net980 net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07714__B _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07206__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06488__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ net575 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06346__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05250__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06100_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[18\] _01782_
+ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07080_ _01619_ _02209_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__nor2_2
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06031_ net157 _01720_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05249__X _00962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06081__A _01762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05215__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06412__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout107 _01650_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_4
XANTENNA__10361__SET_B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout118 net119 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_4
Xfanout129 _01594_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_8
X_07982_ _03319_ _03480_ _03536_ _03535_ _03493_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__o32a_1
X_09721_ _04761_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__inv_2
X_06933_ _02479_ _02485_ _02553_ _02557_ _02603_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a311o_1
XANTENNA__07905__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09652_ _01764_ _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__nor2_1
X_06864_ _02475_ _02494_ _02530_ _02534_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_2_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08603_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01197_ net243 vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__a21oi_1
X_05815_ _00713_ _01501_ _01504_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__a21o_1
X_09583_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ _04665_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__and3_1
X_06795_ _00695_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1
+ vccd1 vccd1 _02466_ sky130_fd_sc_hd__and2_1
XANTENNA__06191__A2 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ _03967_ _03974_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05746_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[8\] _00771_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] vssd1 vssd1 vccd1 vccd1
+ _01446_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_78_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07640__A _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06479__B1 _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ net419 _00676_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__o21a_1
X_05677_ net445 _01297_ _01372_ _01388_ net442 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07416_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\] _03003_
+ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08396_ net459 _03870_ _03843_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_34_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07691__A2 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06256__A _00684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07347_ net415 _00711_ _00796_ _01175_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row
+ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__o41a_1
XFILLER_0_66_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07278_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09017_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ _04274_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05454__A1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06651__B1 _02178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06229_ _01888_ _01898_ _01908_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[1\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold150 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10188__RESET_B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[15\] vssd1 vssd1
+ vccd1 vccd1 net831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[21\] vssd1 vssd1
+ vccd1 vccd1 net853 sky130_fd_sc_hd__dlygate4sd3_1
X_10835__511 vssd1 vssd1 vccd1 vccd1 _10835__511/HI net511 sky130_fd_sc_hd__conb_1
Xhold194 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[14\] vssd1 vssd1
+ vccd1 vccd1 net864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06954__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07815__A _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09919_ net845 net154 net152 _04899_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__a22o_1
XANTENNA__06706__A1 _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05989__B _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09408__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05070__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10625_ clknet_leaf_49_wb_clk_i _00489_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10556_ clknet_leaf_19_wb_clk_i _00424_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10487_ clknet_leaf_23_wb_clk_i _00355_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07198__A1 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05245__A _00684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09940__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06173__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05600_ _01307_ _01308_ _01310_ _01312_ vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__o211a_1
X_06580_ net126 _01642_ _01699_ _02230_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a31o_2
XFILLER_0_87_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05920__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05531_ net424 net423 _01231_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ _01206_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07122__B2 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08275__B _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05251__Y _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08250_ _01384_ _03728_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__nand2_1
X_05462_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right _00963_
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up vssd1 vssd1
+ vccd1 vccd1 _01175_ sky130_fd_sc_hd__or4b_4
XFILLER_0_129_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07201_ _02846_ _02849_ _02850_ _02851_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08181_ net474 net473 vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05393_ _01056_ _01063_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_9_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07132_ _01676_ _01678_ net164 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07063_ _01678_ _01903_ _01935_ _02715_ _02717_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a41o_1
XANTENNA__05436__B2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06523__B net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06014_ net197 _01668_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06400__A3 _02073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07965_ _00753_ net109 vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09704_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\] _04749_ vssd1
+ vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__and2_1
X_06916_ _02496_ _02581_ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__or2_1
X_07896_ _01692_ _03378_ _03406_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__a21o_1
X_09635_ _04699_ _04700_ vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06847_ net432 _02508_ net257 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout268_X net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09566_ net414 _01417_ _01476_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__or3_2
X_06778_ net427 _00986_ net201 _00983_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06538__X _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] _03979_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__a21oi_1
X_05729_ net476 _00796_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09497_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] _00667_
+ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07664__A2 _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08861__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ net927 _03921_ _03653_ vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08379_ _03718_ _03853_ _03854_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__nor3_1
X_10410_ clknet_leaf_23_wb_clk_i _00301_ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_78_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10009__Q team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10341_ clknet_leaf_54_wb_clk_i _00281_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08949__A_N net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10272_ clknet_leaf_73_wb_clk_i _00264_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout83_X net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09463__C net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\] vssd1 vssd1
+ vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
Xfanout471 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[2\] vssd1
+ vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_1
Xfanout482 net483 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_2
X_10987__628 vssd1 vssd1 vccd1 vccd1 _10987__628/HI net628 sky130_fd_sc_hd__conb_1
XANTENNA__05065__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_79_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07104__A1 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10608_ clknet_leaf_47_wb_clk_i _00472_ net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10539_ clknet_leaf_21_wb_clk_i _00407_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09935__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06394__A2 _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__A1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04962_ net1111 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
X_07750_ _01083_ net147 vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__nor2_1
XANTENNA__09868__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06701_ _01699_ _02266_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__nand2_1
X_07681_ _03098_ _03099_ _03144_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__and3_1
XANTENNA__07343__A1 _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09420_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\]
+ _04567_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a21o_1
X_06632_ _02268_ _02272_ _02288_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09351_ net226 _04522_ _04523_ net412 net1126 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__a32o_1
X_06563_ _02153_ _02234_ _02235_ _02236_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06518__B _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05514_ net424 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ _01226_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_74_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08302_ team_07_WB.instance_to_wrap.team_07.heartPixel team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\] vssd1 vssd1 vccd1
+ vccd1 _03780_ sky130_fd_sc_hd__nor3_1
X_09282_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__and4_1
XFILLER_0_118_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06494_ _02155_ _02167_ _02153_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__o21a_1
XANTENNA__07646__A2 _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08233_ _03698_ _03711_ net486 vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05445_ _01011_ _01059_ _01083_ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ _03645_ _03647_ vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05376_ net192 _01015_ _01088_ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__o21a_1
XANTENNA__06534__A _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05409__A1 _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07115_ net283 net88 _01635_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08095_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[12\]
+ _00814_ net483 vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload70 clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload70/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07046_ _02138_ net84 _02699_ _02700_ _02362_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_73_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload81 clknet_leaf_47_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_11_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__04989__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08997_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ _04265_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__or4_1
XANTENNA__07582__A1 _02842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ net268 _03414_ _03416_ _00747_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06137__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ _03433_ _03429_ _03426_ _03425_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__o2bb2a_1
X_09618_ _04666_ _04687_ _04689_ _04664_ net1030 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__a32o_1
X_10890_ net647 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_66_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09549_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[43\]
+ net273 net293 net224 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07098__B1 _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10324_ clknet_leaf_54_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[1\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10255_ clknet_leaf_73_wb_clk_i _00247_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10186_ clknet_leaf_82_wb_clk_i net693 net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08770__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07573__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout290 net293 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_2
XFILLER_0_88_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload6_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07722__B net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07876__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06619__A _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06338__B _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07628__A2 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05230_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\] team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__nor2_2
XFILLER_0_115_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08045__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08589__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05161_ _00873_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05092_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_90_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08920_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[0\]
+ _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09553__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ net451 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ net455 vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07564__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _01102_ net112 vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__nand2_1
X_08782_ _01455_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__or2_1
X_05994_ _01654_ _01685_ _01683_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_58_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04945_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] vssd1 vssd1 vccd1 vccd1
+ _00685_ sky130_fd_sc_hd__inv_2
X_07733_ net278 _01055_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout178_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ _02069_ _02872_ _03198_ _02040_ _03083_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__a221o_1
X_09403_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[47\]
+ _00813_ _00815_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06615_ _02274_ _02279_ _02266_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a21o_1
X_07595_ _01675_ _03042_ _01671_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_66_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06248__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09334_ _04313_ net227 _04511_ net408 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__a32o_1
X_06546_ net218 net187 _01665_ _02219_ _01664_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_138_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09265_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ net406 net230 _04463_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__a22o_1
X_06477_ _01699_ _01901_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_62_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ net459 _01380_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel
+ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__a21oi_1
X_05428_ _01135_ _01138_ _01139_ _01140_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__or4b_1
XFILLER_0_133_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09196_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ net333 _04407_ net1033 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__a41o_1
XFILLER_0_44_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06264__A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08147_ _03627_ _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__and2_2
X_05359_ net194 _01004_ _01010_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__nor3_1
XFILLER_0_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08078_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00820_ net414 vssd1 vssd1
+ vccd1 vccd1 _03592_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07029_ _02335_ _02349_ _02683_ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10040_ _00060_ _00638_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold10 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09581__Y _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold43 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07823__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold87 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 _00172_ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10942_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.tft_reset vssd1 vssd1 vccd1
+ vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06439__A _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05343__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05869__B2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10873_ net549 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_85_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06818__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07491__B1 _03041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06294__B2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05252__D_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06461__X _02135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10307_ clknet_leaf_44_wb_clk_i net815 net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_10238_ clknet_leaf_82_wb_clk_i net702 net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06349__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10169_ clknet_leaf_10_wb_clk_i _00179_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07733__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05253__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06400_ net188 _01642_ _02073_ net205 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_44_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07380_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\] _02979_
+ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__or2_1
XANTENNA__08564__A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_942 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06331_ team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[1\] team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[2\]
+ _01962_ _02006_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireHighlightDetect
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09050_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ _04301_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_13_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07482__B1 _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05700__B net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06262_ net458 net159 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_13_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05213_ _00924_ _00925_ _00923_ vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__or3b_1
XFILLER_0_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08001_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__xor2_1
X_06193_ net215 _01670_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold502 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\] vssd1 vssd1
+ vccd1 vccd1 net1172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[34\]
+ vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05144_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09952_ clknet_leaf_55_wb_clk_i _00067_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_05075_ _00670_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] _00801_
+ _00802_ _00800_ vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08903_ _01401_ _01405_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__nor2_1
X_09883_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\] _01773_ vssd1
+ vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__xnor2_1
X_08834_ net988 _04142_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__nand2_1
X_08765_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] net981 net235 vssd1
+ vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05977_ _01657_ net172 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ _03114_ _03271_ _03269_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__a21o_1
X_04928_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1 vssd1
+ vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
XANTENNA__06259__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08696_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _04114_ _04116_ vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07081__C net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07647_ _01645_ net144 _01741_ net255 vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_64_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07578_ net121 _03135_ _03132_ _02096_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__a211o_1
XANTENNA__06546__X _02220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09317_ net229 _04498_ _04500_ net404 net1024 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_81_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06529_ _01712_ _02088_ _02201_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06276__A1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09248_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ _04449_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09179_ net210 _04398_ _04400_ net402 net1082 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__a32o_1
XFILLER_0_121_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07818__A _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06579__A2 _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08973__A0 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XANTENNA__07537__B net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XANTENNA__06441__B net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XANTENNA__05338__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XANTENNA__07528__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ clknet_leaf_42_wb_clk_i _00102_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[14\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07528__B2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06200__A1 _01863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05344__Y _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10925_ net670 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XANTENNA__07700__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10856_ net532 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_67_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10787_ clknet_leaf_12_wb_clk_i _00608_ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_54_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07545__A2_N _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06019__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08964__A0 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05248__A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10852__528 vssd1 vssd1 vccd1 vccd1 _10852__528/HI net528 sky130_fd_sc_hd__conb_1
X_05900_ _01579_ _01581_ _01584_ _01587_ _01593_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a41oi_4
X_06880_ net108 _02550_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__nand2_1
XANTENNA__06727__C1 _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05831_ _00714_ _01509_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08550_ _03611_ _04003_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__nand2_1
X_05762_ _01459_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\] _01460_ vssd1 vssd1
+ vccd1 vccd1 _01461_ sky130_fd_sc_hd__or4bb_2
XTAP_TAPCELL_ROW_85_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07501_ net96 _01631_ _02009_ _00755_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__and4bb_1
X_05693_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[4\] _01398_ _01400_
+ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[5\] vssd1 vssd1 vccd1 vccd1
+ _01406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08481_ net760 _03952_ net130 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07432_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\] _03013_
+ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07363_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[6\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__and4b_1
XFILLER_0_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09102_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ _04342_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06314_ _01989_ _01988_ _01987_ _01986_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__and4b_1
XFILLER_0_115_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07294_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ _02919_ _02923_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[8\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09033_ _04291_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06245_ net280 _01920_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__nand2_2
XFILLER_0_72_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold310 _00028_ vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__dlygate4sd3_1
X_06176_ net175 net117 net110 net185 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold321 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_up vssd1
+ vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05218__C1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05127_ _00835_ _00836_ _00837_ _00839_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__o2bb2a_1
Xhold354 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold365 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 _00020_ vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold387 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\] vssd1 vssd1
+ vccd1 vccd1 net1057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__dlygate4sd3_1
X_05058_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ _00787_ vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__and3_1
X_09935_ net466 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09866_ net1062 net263 _04865_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_107_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _01448_ _04160_ net1036 vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_29_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _04797_ _04810_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07930__B2 _01067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08748_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ net238 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_2_0_wb_clk_i_X clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ _04058_ _04073_ _04100_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10710_ clknet_leaf_71_wb_clk_i _00541_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06497__A1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06717__A _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05621__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10641_ clknet_leaf_45_wb_clk_i _00505_ net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05572__C_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06436__B net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10572_ clknet_leaf_25_wb_clk_i _00440_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08651__B _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08946__B1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_cleared vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06171__B net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05068__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10955__596 vssd1 vssd1 vccd1 vccd1 _10955__596/HI net596 sky130_fd_sc_hd__conb_1
X_10006_ clknet_leaf_42_wb_clk_i _00026_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07921__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06488__A1 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ net574 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_15_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10839_ net515 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_54_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09938__A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05250__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06030_ net156 _01720_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06362__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05215__A2 team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06412__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout108 net110 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08952__A3 _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout119 net120 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_4
X_07981_ _01692_ _03475_ _03473_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09720_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\] _04754_ vssd1 vssd1
+ vccd1 vccd1 _04761_ sky130_fd_sc_hd__and4_1
X_06932_ _02543_ _02554_ _02549_ _02551_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_52_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09651_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__and2_1
XANTENNA__06176__B1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06863_ net115 _02471_ _02531_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07912__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08602_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\] _04034_
+ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__and2_1
X_05814_ _00713_ _01501_ _01504_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__a21oi_1
X_09582_ _04666_ _04664_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05923__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06794_ net90 _02409_ _02413_ _02438_ _02465_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recPLAYER.playerDetect
+ sky130_fd_sc_hd__o311a_1
XANTENNA__07480__X _03041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08533_ _03977_ _03990_ _03991_ _03989_ vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__a31o_1
X_05745_ _01443_ _01445_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[7\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout160_A _01557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout258_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__B _02744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08464_ net462 _03934_ _03935_ net420 _00731_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__o221a_1
XFILLER_0_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05676_ net442 _01323_ vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07415_ _03003_ net233 _03002_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[11\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_135_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08395_ _01253_ _03733_ _03869_ net460 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_34_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06256__B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07346_ _00965_ _02953_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07277_ net752 _02909_ _02912_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[14\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06543__Y _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07368__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09016_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ _04274_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__a21o_1
X_06228_ _01738_ _01743_ _01899_ _01900_ _01907_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08928__A0 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06159_ net186 _01804_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_76_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold140 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__A3 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold151 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.rand_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold162 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataDc vssd1 vssd1
+ vccd1 vccd1 net832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _00324_ vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__dlygate4sd3_1
X_10874__550 vssd1 vssd1 vccd1 vccd1 _10874__550/HI net550 sky130_fd_sc_hd__conb_1
Xhold184 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[15\] vssd1 vssd1
+ vccd1 vccd1 net854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\] vssd1 vssd1
+ vccd1 vccd1 net865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09918_ _01782_ _04898_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__nand2_1
XANTENNA__07815__B _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09849_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\] _04850_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a21o_1
XANTENNA__06706__A2 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05335__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07831__A _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10030__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06447__A _02086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05989__C net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10624_ clknet_leaf_48_wb_clk_i _00488_ net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10555_ clknet_leaf_19_wb_clk_i _00423_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06642__A1 _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10486_ clknet_leaf_23_wb_clk_i _00354_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09344__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output54_A net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05530_ _01197_ _01241_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06357__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07122__A2 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05461_ _01047_ _01173_ _00964_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07200_ _02040_ _02758_ _02836_ _02848_ _02761_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a32o_1
X_08180_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\] _00704_
+ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_31_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05392_ _00669_ net397 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__nand2_2
XFILLER_0_55_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07131_ net137 net105 net164 vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07062_ net121 _01903_ _01935_ _02716_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__and4_1
XANTENNA__06633__A1 _02119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10858__534 vssd1 vssd1 vccd1 vccd1 _10858__534/HI net534 sky130_fd_sc_hd__conb_1
XFILLER_0_3_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06013_ _01641_ _01674_ _01696_ _01705_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[1\]
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_113_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07189__A2 _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08386__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07964_ net136 _03307_ _03487_ _03490_ _03293_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__o311a_1
XFILLER_0_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ net250 _04749_ _04748_ _04733_ vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__a211oi_1
X_06915_ _01651_ _02497_ _02581_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__or3_1
XANTENNA__06149__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07895_ _03448_ _03449_ _03335_ _03440_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__or4bb_1
XANTENNA_fanout375_A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\] _04698_ vssd1
+ vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nand2_1
XANTENNA__05155__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06846_ _02513_ _02516_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09565_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ net764 net240 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout163_X net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06777_ net427 _00985_ net198 _00971_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08516_ net1118 _03979_ vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__xor2_1
X_05728_ net476 _01432_ _01431_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__a21o_1
X_09496_ net968 net208 _04624_ vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__o21a_1
XANTENNA__07113__A2 _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08447_ _03630_ _03906_ _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05659_ _01322_ _01326_ vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08378_ _00711_ _00727_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08074__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07329_ _02943_ _01040_ _00964_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10340_ clknet_leaf_54_wb_clk_i _00280_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_115_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10271_ clknet_leaf_73_wb_clk_i _00263_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09574__B1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07826__A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10338__RESET_B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 team_07_WB.instance_to_wrap.team_07.memGen.stage\[0\] vssd1 vssd1 vccd1
+ vccd1 net450 sky130_fd_sc_hd__buf_2
Xfanout461 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\] vssd1 vssd1
+ vccd1 vccd1 net461 sky130_fd_sc_hd__buf_2
Xfanout472 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[1\] vssd1
+ vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_2
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__buf_2
XANTENNA__05065__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07561__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05081__A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06863__A1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout90 _01606_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10607_ clknet_leaf_48_wb_clk_i _00471_ net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_86_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10538_ clknet_leaf_21_wb_clk_i _00406_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10469_ clknet_leaf_25_wb_clk_i net736 net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_back
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10970__611 vssd1 vssd1 vccd1 vccd1 _10970__611/HI net611 sky130_fd_sc_hd__conb_1
XANTENNA__07591__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04961_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\] vssd1 vssd1
+ vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
X_06700_ _01740_ _02283_ _02372_ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__o21ai_1
X_07680_ net203 _01700_ _01723_ _02829_ _02835_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__o311a_1
XFILLER_0_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06631_ _02109_ _02301_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__nand2_1
X_09350_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ _04520_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__or2_1
X_06562_ _02148_ _02170_ _02176_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10929__579 vssd1 vssd1 vccd1 vccd1 _10929__579/HI net579 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_47_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08301_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05513_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ _01223_ _01201_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__a211o_1
X_09281_ net228 _04473_ _04474_ net401 net1164 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__a32o_1
X_06493_ net131 net124 _01684_ _02061_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__o31a_1
XFILLER_0_118_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09398__A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08232_ net488 _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_99_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05444_ _01023_ _01080_ _01090_ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_34_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06815__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08163_ _03635_ _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_136_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05375_ net193 _01004_ _01014_ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout123_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06534__B _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07114_ _01811_ _02282_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08094_ _03599_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[12\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload60 clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__inv_8
XFILLER_0_42_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07045_ net286 _00757_ _02697_ _02699_ _01920_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a32o_1
Xclkload71 clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload71/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_73_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload82 clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_73_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10431__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07031__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08996_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__or4b_1
XFILLER_0_76_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07947_ _03500_ _03501_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__nand2_1
XANTENNA__09859__A1 _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout280_X net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ _03345_ _03399_ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__and3_1
X_09617_ _04688_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__inv_2
X_06829_ _02498_ _02499_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06542__B1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ net933 net209 _04653_ vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07098__A1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09479_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] _00667_
+ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__or3_1
XFILLER_0_136_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06845__A1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08047__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10323_ clknet_leaf_54_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[0\]
+ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09547__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10254_ clknet_leaf_73_wb_clk_i _00246_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06460__A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10185_ clknet_leaf_86_wb_clk_i net451 net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10101__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07573__A2 _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout280 _00650_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_4
Xfanout291 net293 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__buf_2
XFILLER_0_89_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06533__B1 _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08038__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05160_ _00848_ _00849_ _00854_ _00872_ vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09946__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05091_ net481 _00811_ _00816_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__and3_2
XFILLER_0_40_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10820__496 vssd1 vssd1 vccd1 vccd1 _10820__496/HI net496 sky130_fd_sc_hd__conb_1
XFILLER_0_126_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08061__S net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06370__A net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09002__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ net296 net294 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ _04185_ vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07801_ _01049_ net99 vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__xnor2_1
X_08781_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[18\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] _04141_ vssd1 vssd1
+ vccd1 vccd1 _04142_ sky130_fd_sc_hd__or4_2
X_05993_ net181 net171 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07732_ _03285_ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__nand2b_1
X_04944_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] vssd1 vssd1 vccd1
+ vccd1 _00684_ sky130_fd_sc_hd__inv_2
XANTENNA__10641__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05714__A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07663_ _03212_ _03216_ _03219_ _03220_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__or4b_1
XFILLER_0_133_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09402_ _00813_ _00815_ _02961_ _04555_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__or4_1
X_06614_ _02269_ _02284_ _02285_ _02286_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07594_ _03152_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09333_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06545_ net214 _01655_ _02054_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_X clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout240_A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout338_A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09264_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ _04462_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06476_ net86 _02148_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__nand2_4
XFILLER_0_117_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08215_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] net459
+ _01270_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08029__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05427_ _01071_ _01096_ _01104_ _01070_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__o22a_1
X_09195_ net1148 net404 net211 _04411_ vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout126_X net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08146_ _03631_ _03632_ _03629_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__o21a_1
X_05358_ _00669_ net397 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08077_ net414 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__nor2_1
X_05289_ net193 _01001_ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__nor2_1
X_07028_ net288 _00754_ net83 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold11 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ _04248_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__o21ai_1
Xhold44 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[1\] vssd1
+ vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[2\] vssd1 vssd1
+ vccd1 vccd1 net769 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_dc vssd1 vssd1
+ vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06439__B _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05869__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10872_ net548 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_27_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05997__C _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06455__A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07491__A1 _03045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10353__RESET_B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10306_ clknet_leaf_45_wb_clk_i net791 net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_10237_ clknet_leaf_82_wb_clk_i net713 net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_10168_ clknet_leaf_10_wb_clk_i _00178_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10213__Q team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10099_ clknet_leaf_31_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.buttonHighlightDetect
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.buttonHighlightPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_63_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05253__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06330_ team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[0\] _02004_ _02005_
+ _01998_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__or4b_1
XFILLER_0_128_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07482__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06261_ _00684_ _01574_ _01575_ _01937_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_13_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08000_ _03550_ _03551_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__xnor2_1
X_05212_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00925_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06192_ net187 net176 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__nand2_4
XANTENNA__10094__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold503 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06037__A2 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05143_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\]
+ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__nand2_1
Xhold514 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07196__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ net7 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
X_05074_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1 vccd1 vccd1
+ _00802_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08902_ net1179 _04216_ net264 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09882_ net847 net153 net151 _04876_ vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08833_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\] _04142_
+ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07942__C1 _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] net1004 net238 vssd1
+ vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__mux2_1
X_05976_ net199 _01667_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07715_ _00754_ _01961_ _03113_ _03270_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__o211ai_1
X_04927_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
X_08695_ net263 _01240_ _04115_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout455_A net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06259__B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07646_ _01728_ _02154_ _01874_ net260 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_105_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07577_ net149 _01685_ net105 vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout243_X net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ _04499_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06528_ _01705_ _02039_ _02060_ _02102_ _02200_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08141__A_N net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09247_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ _04449_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06459_ _02131_ _02132_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08129_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[13\]
+ _03615_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__or2_1
XANTENNA__07818__B net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05236__B1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
X_10022_ clknet_leaf_42_wb_clk_i _00101_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[13\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05906__X _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06751__A3 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input16_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ net669 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10855_ net531 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_116_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10786_ clknet_leaf_14_wb_clk_i _00607_ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07216__A1 _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06019__A2 _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07728__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05248__B _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10417__SET_B net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06727__B1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05830_ _01520_ _01523_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05761_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\] vssd1 vssd1 vccd1
+ vccd1 _01460_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_85_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07500_ _02250_ _02673_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08480_ _03947_ _03951_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__nand2_1
X_05692_ net439 _01404_ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07431_ _03013_ net233 _03012_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[17\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_18_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06366__Y _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07362_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09101_ net212 _04341_ _04343_ net399 net830 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__a32o_1
XFILLER_0_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06313_ net218 _01969_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07293_ _02923_ _02924_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09032_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ _04286_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__and3_1
XANTENNA__07478__X _03039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05466__B1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06244_ net280 _01920_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__and2_2
XANTENNA__06382__X _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06823__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold300 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[34\]
+ vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[39\]
+ vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__dlygate4sd3_1
X_06175_ net187 net114 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout203_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05218__B1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold322 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] vssd1 vssd1
+ vccd1 vccd1 net992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold333 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\] vssd1 vssd1
+ vccd1 vccd1 net1003 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08955__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold344 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__dlygate4sd3_1
X_05126_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\]
+ _00838_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__and3_1
Xhold355 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[23\] vssd1 vssd1
+ vccd1 vccd1 net1025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold366 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\] vssd1 vssd1
+ vccd1 vccd1 net1036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold377 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\] vssd1 vssd1 vccd1
+ vccd1 net1047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold388 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\] vssd1 vssd1
+ vccd1 vccd1 net1058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\] vssd1 vssd1
+ vccd1 vccd1 net1069 sky130_fd_sc_hd__dlygate4sd3_1
X_05057_ _00772_ _00784_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__nor2_1
X_09934_ net1079 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05726__X _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input8_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[1\]
+ net242 _04228_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__and3_1
XANTENNA__08102__X _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06718__B1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ net195 _04165_ vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_29_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\] _04815_ vssd1
+ vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__or2_1
X_08747_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ net238 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__mux2_1
X_05959_ _01574_ _01575_ net145 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__a21o_4
XTAP_TAPCELL_ROW_124_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _04080_ _04102_ _04084_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05902__A _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06497__A2 _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ _03181_ _03185_ _03186_ _02734_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10640_ clknet_leaf_45_wb_clk_i _00504_ net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10571_ clknet_leaf_26_wb_clk_i _00439_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05457__B1 _01113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10028__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08946__A1 _00709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05349__A team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05068__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08037__A_N net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06709__B1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ clknet_leaf_41_wb_clk_i _00025_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05355__Y _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07921__A2 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10140__D team_07_WB.instance_to_wrap.team_07.recPLAYER.playerDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10907_ net573 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_15_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07685__A1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06488__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838_ net514 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05250__C team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10769_ clknet_leaf_66_wb_clk_i _00590_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07739__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06362__B net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06412__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout109 net110 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_2
X_07980_ _01679_ _03492_ _03495_ _03534_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__o22a_1
XANTENNA__07474__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06931_ _02543_ _02548_ _02559_ _02471_ net95 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__o32a_1
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09650_ _04713_ _04711_ net1119 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06862_ _02494_ _02532_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__nand2_1
XANTENNA__06176__A1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06176__B2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08601_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared _01239_ vssd1
+ vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05813_ _01492_ _01504_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__xor2_1
X_09581_ _01793_ _03992_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__nor2_2
X_06793_ _02444_ _02456_ _02464_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08532_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\]
+ _03985_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\] vssd1 vssd1
+ vccd1 vccd1 _03991_ sky130_fd_sc_hd__a31o_1
X_05744_ _00766_ _01444_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05722__A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07676__A1 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] net462
+ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__nand2_1
XANTENNA__07676__B2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05675_ _01344_ _01387_ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07414_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\]
+ _02999_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08394_ net461 _03868_ _03840_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07345_ net418 _02953_ _02954_ _00964_ _02955_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing_mod_locator.nxt_mod_col
+ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout320_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07276_ _02912_ _02913_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[13\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06553__A _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09015_ net251 _04277_ _04278_ net403 net1100 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__a32o_1
XFILLER_0_130_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06227_ _01838_ _01902_ _01905_ _01906_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__or4_1
Xhold130 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06158_ _01835_ _01836_ _01838_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__or3_1
Xhold141 _00327_ vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold152 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[6\] vssd1 vssd1
+ vccd1 vccd1 net822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[15\]
+ vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__dlygate4sd3_1
X_05109_ net1049 _00817_ _00823_ net1011 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__a22o_1
Xhold174 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[8\] vssd1 vssd1
+ vccd1 vccd1 net844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[9\] vssd1 vssd1
+ vccd1 vccd1 net855 sky130_fd_sc_hd__dlygate4sd3_1
X_06089_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\] vssd1 vssd1 vccd1
+ vccd1 _01772_ sky130_fd_sc_hd__or3_1
Xhold196 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07384__A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09917_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\] _01781_
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[17\] vssd1 vssd1 vccd1
+ vccd1 _04898_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09848_ net269 _04852_ _04853_ net247 net1174 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__a32o_1
XFILLER_0_77_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] _04803_ vssd1
+ vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_122_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07831__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07116__B1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07323__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07667__B2 _03095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05351__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10623_ clknet_leaf_48_wb_clk_i _00487_ net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ clknet_leaf_20_wb_clk_i _00422_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06642__A2 _02209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10485_ clknet_leaf_13_wb_clk_i _00353_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09041__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07658__A1 _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08855__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05460_ _00968_ _01166_ _01172_ _01162_ _01165_ vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05391_ net435 _00967_ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07130_ _01694_ net164 _02775_ _02767_ _02762_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__a32o_1
XFILLER_0_55_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06373__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07061_ _01639_ _02714_ _02335_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_97_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06012_ _01704_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07963_ _03398_ _03401_ _03516_ _03517_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_71_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09702_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[8\] _04742_ vssd1 vssd1
+ vccd1 vccd1 _04749_ sky130_fd_sc_hd__and4_1
X_06914_ _02535_ _02584_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__nand2_1
XANTENNA__06149__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07894_ net106 _01692_ net186 vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09633_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\] _04698_ vssd1
+ vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__or2_1
X_06845_ net201 _02500_ _02515_ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout368_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ net776 net236 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__mux2_1
X_06776_ _00984_ net174 _02447_ net183 vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__o22a_1
XFILLER_0_136_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08515_ _00698_ _03976_ _03979_ vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__a21oi_1
X_05727_ _01432_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__inv_2
X_09495_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[19\]
+ net272 _04623_ net290 net221 vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout156_X net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08446_ _03908_ _03919_ net490 _03753_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05658_ _01255_ _01278_ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08377_ _03835_ _03852_ net489 vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05589_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\] vssd1 vssd1 vccd1
+ vccd1 _01302_ sky130_fd_sc_hd__or3b_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07328_ _02942_ _02419_ _01109_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07259_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[8\]
+ _02900_ _02902_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[8\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09023__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ clknet_leaf_73_wb_clk_i _00262_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07585__B1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout440 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[1\] vssd1 vssd1 vccd1
+ vccd1 net440 sky130_fd_sc_hd__buf_2
Xfanout451 net452 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_2
XANTENNA__05346__B _01000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout462 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\] vssd1 vssd1
+ vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_2
Xfanout473 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[1\] vssd1
+ vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout484 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07561__B _02744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06458__A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06560__A1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06177__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08225__A_N net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924__669 vssd1 vssd1 vccd1 vccd1 net669 _10924__669/LO sky130_fd_sc_hd__conb_1
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06464__Y _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout91 net92 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__buf_2
XFILLER_0_80_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_88_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10606_ clknet_leaf_48_wb_clk_i _00470_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10537_ clknet_leaf_20_wb_clk_i _00405_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_17_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10468_ clknet_leaf_20_wb_clk_i net739 net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_select
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07736__B _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10399_ clknet_leaf_10_wb_clk_i net673 net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07591__A3 _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04960_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\] vssd1 vssd1
+ vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06630_ _02291_ _02299_ _02302_ _02259_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a31o_1
XANTENNA__06551__A1 _02220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06561_ _02067_ _02150_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__nor2_2
XFILLER_0_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08300_ _03777_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05512_ net424 _01221_ _01222_ _01224_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__a22o_1
X_09280_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__nand3_1
X_10825__501 vssd1 vssd1 vccd1 vccd1 _10825__501/HI net501 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_47_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06492_ _02076_ _02155_ _02153_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08231_ _03708_ _03709_ _03702_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__o21a_1
X_05443_ _01061_ _01070_ _01094_ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06374__Y _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06815__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08162_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[3\] _03639_
+ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__nand2_1
XANTENNA__08056__A1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05374_ net194 _01013_ _01086_ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__o21a_1
XANTENNA__08056__B2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07113_ _01634_ _02332_ _02766_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08093_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[11\]
+ _00814_ net483 vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout116_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload50 clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_30_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07044_ _02088_ _02698_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__nor2_2
Xclkload61 clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__inv_6
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload72 clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__inv_6
XANTENNA__06831__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload83 clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06550__B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07031__A2 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05166__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07946_ net275 _03414_ _03416_ _00752_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__o22ai_1
XANTENNA__09859__A2 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07662__A _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07877_ _01145_ net112 _03431_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout273_X net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\] _04682_ vssd1 vssd1
+ vccd1 vccd1 _04688_ sky130_fd_sc_hd__and4_1
X_06828_ net432 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1 vssd1
+ vccd1 vccd1 _02499_ sky130_fd_sc_hd__nor2_1
XANTENNA__06542__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05182__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06759_ net219 _02419_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__nand2_1
X_09547_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[42\]
+ net273 net293 net224 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09478_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[15\]
+ net222 _04605_ net923 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10231__SET_B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08429_ _03639_ _03899_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__o21a_1
XANTENNA__05648__A3 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06284__Y _01961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08047__A1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload0 clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_18_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10993__634 vssd1 vssd1 vccd1 vccd1 _10993__634/HI net634 sky130_fd_sc_hd__conb_1
X_10322_ clknet_leaf_44_wb_clk_i net750 net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_10253_ clknet_leaf_73_wb_clk_i _00245_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06460__B _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07558__B1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ clknet_leaf_86_wb_clk_i net454 net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07573__A3 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout270 net271 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_2
XANTENNA__07572__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout281 _00650_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_2
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08955__X _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08038__A1 _00706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06049__B1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05090_ _00813_ _00815_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06370__B _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07800_ _01078_ net94 vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__xnor2_1
X_08780_ net411 _01453_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05992_ net181 net171 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__nor2_2
XANTENNA__06772__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06772__B2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07731_ _01105_ net276 _01625_ _01636_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__a31o_1
X_04943_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\] vssd1
+ vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
XANTENNA__05980__C1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07662_ _01904_ _02765_ _03071_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__or3_1
XANTENNA__05714__B _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09401_ _02962_ _03592_ _04556_ _02963_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__o2bb2a_1
X_06613_ _01653_ _02270_ net254 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07593_ _01610_ _02298_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__nand2_2
XANTENNA__05878__A3 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09332_ net227 net411 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__mux2_1
X_06544_ net97 _02131_ _02215_ _02217_ _02211_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a41o_1
XFILLER_0_133_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09263_ net230 _04461_ _04462_ net406 net1171 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06475_ net86 _02148_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__and2_2
X_08214_ _01293_ _03676_ _03692_ net460 vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__o22a_1
XANTENNA__08029__A1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05426_ _00966_ _01081_ _01050_ _01036_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__a2bb2o_1
X_09194_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__xnor2_1
X_10977__618 vssd1 vssd1 vccd1 vccd1 _10977__618/HI net618 sky130_fd_sc_hd__conb_1
XFILLER_0_105_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08145_ net467 net470 vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__nor2_1
X_05357_ net191 _01005_ _01021_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout400_A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout119_X net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08076_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ net395 net297 net981 _03590_ vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__a221o_1
X_05288_ _00996_ _01000_ vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__or2_1
XANTENNA__06561__A _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07027_ _02677_ _02681_ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09872__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold12 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__o21a_1
Xhold45 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _01078_ net200 _03312_ _01068_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__o22a_1
Xhold78 _00116_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__dlygate4sd3_1
X_10940_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sdi vssd1 vssd1
+ vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06515__A1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05318__A2 _01014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10871_ net547 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_79_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09465__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_9 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07567__A _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10305_ clknet_leaf_45_wb_clk_i _00043_ net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10236_ clknet_leaf_76_wb_clk_i net718 net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_10167_ clknet_leaf_7_wb_clk_i _00177_ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_89_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10098_ clknet_leaf_80_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[3\]
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.labelPixel\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07703__B1 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06260_ _01677_ _01936_ net458 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__mux2_1
XANTENNA__07482__A2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10339__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05211_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00924_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_13_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06191_ net218 net101 net91 net199 _01871_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05142_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\]
+ vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__nand2_1
Xhold504 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\] vssd1 vssd1
+ vccd1 vccd1 net1174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08072__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06381__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07196__B _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05073_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1 vccd1 vccd1
+ _00801_ sky130_fd_sc_hd__nand2_1
X_09950_ net464 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08901_ _01404_ _04198_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09881_ _01773_ _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08832_ _04142_ _04175_ net196 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07942__B1 _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05725__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08763_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ net235 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__mux2_1
X_05975_ net260 net172 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_68_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout183_A _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07714_ net97 _02217_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04926_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\] vssd1
+ vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
X_08694_ _04112_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__nand2_2
XFILLER_0_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07645_ _03180_ _03187_ _03191_ _03202_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__or4b_1
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07576_ net141 net169 net164 net137 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09315_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04494_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06527_ net135 _01698_ _02056_ _02091_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__or4_1
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout236_X net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09246_ net230 _04448_ _04450_ net407 net871 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__a32o_1
X_06458_ net205 _02112_ _02113_ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__or3_1
XFILLER_0_134_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05409_ _01083_ _01087_ _01093_ _01098_ _01082_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_16_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09177_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ _04396_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__and2_1
XANTENNA__06681__B1 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06389_ _02060_ _02061_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08128_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[12\]
+ _03614_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08059_ net454 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ net393 net296 vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XANTENNA_fanout96_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_0_101_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XANTENNA__07460__A_N net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
X_10021_ clknet_leaf_42_wb_clk_i _00100_ net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[12\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_129_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05922__X _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07850__A _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923_ net668 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
XFILLER_0_86_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07700__A3 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10854_ net530 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__06466__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ clknet_leaf_66_wb_clk_i _00606_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.audio
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06672__B1 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07216__A2 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06019__A3 _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05248__C _00960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10224__Q team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10781__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10219_ clknet_leaf_90_wb_clk_i _00223_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07924__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09677__A0 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05760_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\] _01458_
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[4\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_85_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05691_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\] _00796_
+ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__nand2_1
XANTENNA__07152__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07430_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\]
+ _03009_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06376__A _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07361_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06312_ net200 _01966_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09100_ _04342_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07292_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06663__X _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09031_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ _04286_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06243_ net283 net277 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__nor2_1
XANTENNA__07928__A1_N _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06174_ net215 net96 net94 net197 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a22o_1
Xhold301 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[6\] vssd1 vssd1 vccd1
+ vccd1 net971 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold312 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[1\] vssd1 vssd1
+ vccd1 vccd1 net982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[38\]
+ vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__dlygate4sd3_1
X_05125_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__nand2_1
XANTENNA__08955__A2 _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\] vssd1 vssd1
+ vccd1 vccd1 net1026 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold367 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\] vssd1 vssd1 vccd1
+ vccd1 net1048 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__dlygate4sd3_1
X_05056_ net1020 _00774_ _00784_ _00786_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[5\]
+ sky130_fd_sc_hd__o31ai_1
X_09933_ net1104 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout398_A _00943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09864_ net860 net263 _04864_ vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__a21o_1
XANTENNA__06718__B2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08815_ net942 _04164_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_107_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _04811_ _04814_ _04816_ _04808_ net1156 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_29_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06194__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout186_X net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08746_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ net238 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__mux2_1
X_05958_ net145 net136 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_124_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04909_ net282 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
XANTENNA__07143__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08677_ _04089_ _04092_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__nor2_1
X_05889_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] _01579_
+ _01581_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07628_ _01660_ _02061_ _03183_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__a21bo_1
XANTENNA__05902__B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07559_ _02135_ _02140_ _02150_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ clknet_leaf_26_wb_clk_i _00438_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04435_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05349__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout99_X net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06709__A1 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ clknet_leaf_42_wb_clk_i _00024_ net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05365__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05067__D_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06908__B _01557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10906_ net572 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XANTENNA__07685__A2 _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06196__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10837_ net513 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_7_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10768_ clknet_leaf_62_wb_clk_i _00589_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05448__A1 _01104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10699_ clknet_leaf_70_wb_clk_i _00530_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06362__C _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06930_ _02533_ _02585_ _02600_ _02569_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a211o_1
XANTENNA__09898__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06861_ _02530_ _02531_ _02475_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06176__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ _03623_ net767 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__o21a_1
X_05812_ _01492_ _01504_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__xnor2_1
X_09580_ _01793_ _03967_ _03976_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__o21ai_2
X_06792_ net113 _02458_ _02463_ _02457_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08531_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\] _03985_ vssd1 vssd1
+ vccd1 vccd1 _03990_ sky130_fd_sc_hd__nand4_1
X_05743_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\]
+ _00775_ _00652_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07852__A1_N net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05674_ net421 _01258_ _01381_ _01386_ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__a211o_1
X_08462_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] _03686_
+ _03688_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07676__A2 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07413_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\]
+ _02998_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\] vssd1
+ vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__a31o_1
X_08393_ _01257_ _03728_ _03867_ net462 vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07489__X _03050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07344_ net490 net418 vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07275_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09014_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ _04274_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__or2_1
X_06226_ net97 _01878_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08389__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold120 _00105_ vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__dlygate4sd3_1
X_06157_ net96 _01831_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold131 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[1\]
+ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout101_X net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold142 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold153 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__dlygate4sd3_1
X_05108_ net1045 _00817_ _00823_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__a22o_1
Xhold164 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold175 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[17\] vssd1 vssd1
+ vccd1 vccd1 net845 sky130_fd_sc_hd__dlygate4sd3_1
X_06088_ _00654_ _01771_ _01411_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__a21oi_1
Xhold186 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.rand_num\[2\]
+ vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05611__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09916_ net1106 net153 net151 _04897_ vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05039_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__nand4_1
XANTENNA__05185__A team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09847_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\] _04850_ vssd1
+ vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09778_ _04799_ _04800_ _04801_ _04802_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_122_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ net1138 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ net234 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__mux2_1
XANTENNA__07116__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10842__518 vssd1 vssd1 vccd1 vccd1 _10842__518/HI net518 sky130_fd_sc_hd__conb_1
XFILLER_0_64_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10622_ clknet_leaf_48_wb_clk_i _00486_ net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06744__A team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10166__RESET_B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10553_ clknet_leaf_20_wb_clk_i _00421_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10484_ clknet_leaf_13_wb_clk_i _00352_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06478__X _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07107__A1 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07107__B2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07658__A2 _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05390_ net192 _01013_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07060_ _01639_ _02713_ _02714_ _02686_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__o31a_1
XFILLER_0_70_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06011_ net126 _01683_ _01703_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07485__A _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07043__B1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07962_ net262 _01621_ _03392_ _03427_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_71_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09701_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[8\] _04745_ vssd1
+ vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__nor2_1
X_06913_ _00751_ _02486_ _02539_ _02537_ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06149__A2 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07893_ _03306_ _03446_ _03447_ _03445_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__or4b_1
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ _04697_ _04698_ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__nor2_1
X_06844_ net217 _02511_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__nand2_1
X_09563_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ net803 net236 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06775_ _02446_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout263_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] _00657_ _01793_
+ _03977_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__a31o_1
X_05726_ _01108_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back vssd1
+ vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__or3b_4
X_09494_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ _00667_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06267__C net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08445_ net465 _03713_ _03918_ _03911_ net415 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__a311o_1
XFILLER_0_136_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05657_ _01278_ _01369_ vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_93_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10945__586 vssd1 vssd1 vccd1 vccd1 _10945__586/HI net586 sky130_fd_sc_hd__conb_1
XANTENNA_fanout149_X net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08376_ net487 _03846_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__or3_1
X_05588_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07327_ net426 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__mux2_1
XANTENNA__08074__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07258_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[9\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06209_ net91 _01800_ _01824_ _01600_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a22o_1
X_07189_ _01717_ _01737_ _01828_ net202 vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07585__A1 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_2
Xfanout441 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[0\] vssd1 vssd1 vccd1
+ vccd1 net441 sky130_fd_sc_hd__clkbuf_4
Xfanout452 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_4
Xfanout463 net466 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_4
Xfanout474 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[0\] vssd1
+ vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_2
XANTENNA__08938__B _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout485 net487 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06739__A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07334__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06560__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout81 net82 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_2
Xfanout92 _01606_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_2
X_10605_ clknet_leaf_47_wb_clk_i _00469_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10536_ clknet_leaf_21_wb_clk_i _00404_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ clknet_leaf_20_wb_clk_i net731 net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_right
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06480__Y _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06921__B net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07025__B1 _00943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08773__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07576__A1 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06379__A2 _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10398_ clknet_leaf_10_wb_clk_i net724 net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07576__B2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11019_ net643 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_0_95_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06000__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06001__X _01694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06368__B _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06560_ _01739_ net166 _02092_ _02155_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a211o_1
XANTENNA__08864__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05511_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ _01198_ _01203_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__a22o_1
X_10864__540 vssd1 vssd1 vccd1 vccd1 _10864__540/HI net540 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_47_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06491_ net281 net284 net267 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_47_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ _00683_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__nand2_2
X_05442_ _01038_ _01079_ _01067_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_99_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08161_ net475 _03634_ _03639_ net469 vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__a31o_1
X_05373_ _01085_ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07112_ _02332_ net82 _02735_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08092_ net953 _03594_ _03595_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload40 clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__inv_8
XFILLER_0_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07043_ _01675_ _01828_ net203 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload51 clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload51/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload62 clknet_leaf_71_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__inv_8
XFILLER_0_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload73 clknet_leaf_57_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_73_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout109_A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload84 clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__inv_16
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08994_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ _04260_ _04262_ _04258_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__o31a_1
XFILLER_0_76_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07945_ _03480_ _03486_ _03493_ _03499_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__a22o_1
X_07876_ _00970_ net118 net112 _01145_ _03430_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__o221a_1
X_09615_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\]
+ _04682_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\] vssd1 vssd1
+ vccd1 vccd1 _04687_ sky130_fd_sc_hd__a31o_1
X_06827_ net432 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1 vssd1
+ vccd1 vccd1 _02498_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout266_X net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06542__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09546_ net907 net209 _04652_ vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__o21a_1
X_06758_ _02428_ _02429_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_66_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05709_ _01421_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__inv_2
X_09477_ net923 net207 _04611_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__o21a_1
X_06689_ net98 net89 net86 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08428_ _03662_ _03891_ _00703_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload1 clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_22_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08359_ team_07_WB.instance_to_wrap.team_07.borderGen.borderPixel _03719_ _03834_
+ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10321_ clknet_leaf_47_wb_clk_i net788 net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07329__S _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09547__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10252_ clknet_leaf_26_wb_clk_i _00244_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.internalSck
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07558__A1 _01921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05357__B _01005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ clknet_leaf_9_wb_clk_i _00193_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input39_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_4
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_4
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_2
XANTENNA__07572__B net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout293 _04584_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10848__524 vssd1 vssd1 vccd1 vccd1 _10848__524/HI net524 sky130_fd_sc_hd__conb_1
XFILLER_0_69_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08684__A team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07494__B1 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06049__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10519_ clknet_leaf_17_wb_clk_i _00387_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05548__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10935__585 vssd1 vssd1 vccd1 vccd1 _10935__585/HI net585 sky130_fd_sc_hd__conb_1
X_05991_ net214 net184 _01663_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__a21o_2
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07730_ net109 _03280_ _03284_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__or3b_2
XFILLER_0_46_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04942_ net1182 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
XANTENNA__05980__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07661_ _02829_ _03213_ _03218_ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09400_ _02959_ _02961_ _02964_ team_07_WB.instance_to_wrap.ssdec_ss _04556_ vssd1
+ vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__a221o_1
X_06612_ _01720_ _02021_ _02271_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__o21a_1
X_07592_ _01664_ _01669_ _03149_ _03150_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09331_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ net6 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ _04509_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_66_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06543_ net89 _02216_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__nand2_2
XFILLER_0_8_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09262_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ _04459_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_138_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06474_ _01596_ _01603_ _01598_ _01590_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__o211a_4
XFILLER_0_28_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08213_ _01281_ _03679_ _03691_ net461 vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_106_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05425_ net435 _01099_ _01113_ _01085_ _01137_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09193_ net211 _04409_ _04410_ net404 net1165 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__a32o_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08144_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__nand2_2
X_05356_ _00967_ _01062_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__or2_2
XANTENNA__08434__C1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08075_ net454 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__and2b_1
X_05287_ _00675_ _00999_ vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_112_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06561__B _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07026_ _02678_ _02680_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__nor2_1
XANTENNA__08215__A_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] net836
+ net447 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__mux2_1
Xhold24 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[2\]
+ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _01068_ _03312_ net190 _01091_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__a2bb2o_1
Xhold68 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[18\] vssd1 vssd1
+ vccd1 vccd1 net738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[24\] vssd1 vssd1
+ vccd1 vccd1 net749 sky130_fd_sc_hd__dlygate4sd3_1
X_07859_ _03299_ _03413_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__or2_1
X_10870_ net546 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_85_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09529_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[33\]
+ net270 _04643_ net291 net223 vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a221o_1
X_10960__601 vssd1 vssd1 vccd1 vccd1 _10960__601/HI net601 sky130_fd_sc_hd__conb_1
XFILLER_0_137_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06279__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08976__A0 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06451__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10304_ clknet_leaf_47_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[17\]
+ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10235_ clknet_leaf_82_wb_clk_i net712 net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[5\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06203__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06203__B2 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10166_ clknet_leaf_6_wb_clk_i _00176_ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_10097_ clknet_leaf_81_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[2\]
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.labelPixel\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06199__A _01681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10889__646 vssd1 vssd1 vccd1 vccd1 net646 _10889__646/LO sky130_fd_sc_hd__conb_1
XANTENNA__10362__RESET_B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__B2 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload4_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10999_ net637 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_44_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07482__A3 _01901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05210_ _00919_ _00920_ _00921_ _00922_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_13_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07219__B1 _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06190_ net187 net114 _01866_ _01870_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_72_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06662__A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05141_ _00850_ _00851_ _00852_ _00853_ vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__a22o_1
Xhold505 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__dlygate4sd3_1
X_05072_ net427 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1 vssd1
+ vccd1 vccd1 _00800_ sky130_fd_sc_hd__xor2_1
XANTENNA__07196__C _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08900_ _04215_ net903 _04209_ vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__mux2_1
X_09880_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[3\] _01772_ vssd1
+ vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__nand2_1
X_08831_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\]
+ _04141_ net868 vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__o31ai_1
XANTENNA__06745__A2 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__A1 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__B2 _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08762_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__mux2_1
XANTENNA__05725__B net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05974_ net184 net176 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__or2_1
X_07713_ _03256_ _03258_ _03268_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_68_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04925_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] vssd1
+ vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
X_08693_ net243 _04113_ _04040_ _01759_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout176_A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07644_ _03074_ _03192_ _03195_ _03201_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_105_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07575_ _01686_ _02263_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout343_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09314_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ _04491_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__a31o_1
X_06526_ _01687_ _01690_ _02047_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09245_ _04449_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__inv_2
X_06457_ _01711_ _02089_ _02050_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout131_X net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05408_ _01111_ _01112_ _01119_ _01120_ _01073_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__o2111a_1
X_09176_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ _04396_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__or2_1
X_06388_ _02061_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08958__B1 _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08127_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[11\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[10\] _03613_
+ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05339_ net193 _01004_ _01005_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__nor3_2
XFILLER_0_4_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08058_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ net294 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
X_07009_ _02661_ _02665_ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XFILLER_0_101_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10020_ clknet_leaf_42_wb_clk_i net954 net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout89_A _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05916__A _01582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10922_ net667 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
XANTENNA__07850__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07697__B1 _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10853_ net529 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10784_ clknet_leaf_65_wb_clk_i _00605_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10218_ clknet_leaf_86_wb_clk_i _00222_ net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05545__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ clknet_leaf_1_wb_clk_i net719 net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05690_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\] _00796_
+ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10306__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07360_ _02968_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_sck_fl_enable
+ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06311_ net199 _01966_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06521__A2_N _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07291_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ _02922_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__a31o_1
X_09030_ net252 _04288_ _04289_ net407 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__a32o_1
XFILLER_0_127_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06242_ _01827_ _01847_ _01918_ _01919_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[3\]
+ sky130_fd_sc_hd__and4_1
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06392__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06173_ net215 net96 _01853_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a21oi_1
Xhold302 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] vssd1 vssd1
+ vccd1 vccd1 net972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold313 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] vssd1 vssd1
+ vccd1 vccd1 net983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold324 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__dlygate4sd3_1
X_05124_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\]
+ _00835_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__a21o_1
Xhold335 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\] vssd1 vssd1
+ vccd1 vccd1 net1005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold346 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[8\] vssd1
+ vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold357 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\] vssd1 vssd1 vccd1
+ vccd1 net1027 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ net411 _01787_ net892 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__o21a_1
X_05055_ _00766_ _00774_ _00785_ net1020 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__o211ai_1
Xhold368 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\] vssd1 vssd1
+ vccd1 vccd1 net1038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold379 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04911__Y _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10284__RESET_B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09863_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ net241 _04228_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__and3_1
XANTENNA__06179__B1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout293_A _04584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07915__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08814_ _04163_ _04164_ net195 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__a21oi_1
X_09794_ _04815_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07951__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08745_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[19\]
+ net239 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__mux2_1
X_05957_ net132 net125 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__nand2_8
XTAP_TAPCELL_ROW_124_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout179_X net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04908_ net287 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
X_08676_ _04099_ _04101_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__a21o_1
X_05888_ _01578_ _01580_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__nor2_2
XFILLER_0_95_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07627_ _02171_ _03184_ _03183_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07558_ _01921_ _02214_ _01618_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06509_ _00750_ _01611_ _02042_ _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__or4_1
XFILLER_0_134_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07489_ _01730_ _02082_ _03048_ _03049_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09228_ net231 _04436_ _04437_ net408 net872 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09159_ net210 _04385_ _04386_ net401 net883 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__a32o_1
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08946__A3 _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07845__B net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10003_ clknet_leaf_40_wb_clk_i _00023_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input21_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07861__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06477__A _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05381__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10905_ net571 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_54_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10836_ net512 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08095__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10767_ clknet_leaf_62_wb_clk_i _00588_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06645__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06645__B2 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10698_ clknet_leaf_70_wb_clk_i _00529_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07755__B net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06860_ net90 _02474_ _02529_ net108 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_52_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05811_ _00713_ _01492_ net219 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__or3_1
X_06791_ net113 _02458_ _02462_ net118 _02461_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08530_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\] _03978_ vssd1
+ vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__and2_1
X_05742_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\] _00775_ _00783_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\] vssd1 vssd1 vccd1 vccd1
+ _01443_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08322__A1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08461_ net822 net130 _03933_ vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__o21ba_1
X_05673_ _01276_ _01279_ _01300_ _01385_ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__a31o_1
X_07412_ net992 _02999_ _03001_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[10\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08392_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08086__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07450__A_N net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07343_ _01109_ _02953_ _00710_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06393__Y _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout139_A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09210__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07274_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ _01389_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09013_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ _04274_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06225_ _01812_ _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout306_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold110 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__dlygate4sd3_1
X_06156_ net91 _01834_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__nand2_1
Xhold121 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 _00166_ vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold143 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__dlygate4sd3_1
X_05107_ net481 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ _00821_ _00817_ net1015 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__a32o_1
XANTENNA__07061__A1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold154 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__dlygate4sd3_1
X_06087_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] _01771_ _01411_
+ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a21o_1
Xhold176 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 team_07_WB.instance_to_wrap.ssdec_sck vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold198 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[18\] vssd1 vssd1
+ vccd1 vccd1 net868 sky130_fd_sc_hd__dlygate4sd3_1
X_05038_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[13\]
+ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__and4b_1
X_09915_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\] _01781_
+ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05185__B team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\] _04850_ vssd1
+ vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08561__A1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07681__A _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09777_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[14\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__or4bb_1
X_06989_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\]
+ _02651_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\] vssd1
+ vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__a31o_1
XANTENNA__06572__B1 _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08728_ net1043 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05913__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07116__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08659_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ _04049_ _04051_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06324__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06584__X team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10881__557 vssd1 vssd1 vccd1 vccd1 _10881__557/HI net557 sky130_fd_sc_hd__conb_1
XFILLER_0_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10621_ clknet_leaf_48_wb_clk_i _00485_ net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10771__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10552_ clknet_leaf_20_wb_clk_i _00420_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10483_ clknet_leaf_22_wb_clk_i _00351_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05928__X _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10135__RESET_B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06563__B1 _02235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05382__Y _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05823__B _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06866__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08068__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ net495 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_138_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06618__A1 _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06618__B2 _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06010_ net135 net170 net141 _01683_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07043__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07485__B _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07961_ _01689_ _03380_ _03388_ _01679_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__o22a_1
X_09700_ _04734_ _04746_ _04747_ vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06912_ net107 _02493_ _02575_ _02582_ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__or4_1
X_07892_ _01091_ net178 vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__xor2_1
X_09631_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\]
+ _04696_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06843_ net201 _02500_ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05292__Y _01005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ net779 net240 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__mux2_1
X_06774_ net426 _00973_ _00985_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08513_ _00698_ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__nor2_1
X_05725_ net476 net491 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09493_ net929 net208 _04622_ vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout256_A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08444_ net485 _03881_ _03917_ _03722_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__o31ai_1
X_05656_ _01280_ _01331_ _01337_ _01342_ _01368_ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__a41o_1
XFILLER_0_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08375_ _03709_ _03848_ _03850_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__o21a_1
X_05587_ _01295_ _01299_ vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07326_ _02939_ _02941_ _02936_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[1\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07257_ _02898_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[7\]
+ _02901_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[7\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06208_ _01837_ _01845_ _01835_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07188_ _02277_ _02836_ _02829_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06139_ _01809_ _01817_ _01818_ _01819_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07346__A_N _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07585__A2 _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout420 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] vssd1
+ vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout431 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_4
Xfanout442 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[2\] vssd1 vssd1 vccd1
+ vccd1 net442 sky130_fd_sc_hd__buf_2
Xfanout453 net455 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_2
Xfanout464 net465 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_2
Xfanout475 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[0\] vssd1
+ vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05924__A _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout486 net487 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_2
X_09829_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\] _04838_ vssd1
+ vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__and2_1
XANTENNA__06545__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08300__A _03777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06739__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11024__644 vssd1 vssd1 vccd1 vccd1 _11024__644/HI net644 sky130_fd_sc_hd__conb_1
XFILLER_0_138_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05520__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05520__B2 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10604_ clknet_leaf_47_wb_clk_i _00468_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout82 _02731_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout93 net94 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_4
XFILLER_0_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10535_ clknet_leaf_21_wb_clk_i _00403_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10466_ clknet_leaf_20_wb_clk_i net732 net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_left
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06490__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07025__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10397_ clknet_leaf_10_wb_clk_i net882 net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07576__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06379__A3 _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11018_ net391 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_26_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06000__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08864__B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05510_ net424 net422 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__nand2b_2
X_06490_ net287 net279 _00748_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__and3_4
XFILLER_0_28_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05441_ _01030_ _01097_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08160_ net471 _03644_ _03634_ vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__mux2_1
X_05372_ net191 _01014_ _01019_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__nor3_1
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10905__571 vssd1 vssd1 vccd1 vccd1 _10905__571/HI net571 sky130_fd_sc_hd__conb_1
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07111_ _02764_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08091_ _03598_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[10\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload30 clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_6
Xclkload41 clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__inv_6
X_07042_ _02086_ _02696_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__and2_2
Xclkload52 clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload63 clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__inv_8
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload74 clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_73_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload85 clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__05287__Y _01000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08993_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04261_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_110_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10423__Q team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07944_ _03496_ _03498_ _03495_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07875_ _00970_ net118 _03349_ _03423_ _03348_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09614_ _04685_ _04686_ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__nand2_1
X_06826_ _02495_ _02496_ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__nand2_1
X_09545_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[41\]
+ net273 net293 net225 vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__a211o_1
X_06757_ net257 _02427_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout161_X net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05708_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _01419_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__or3_2
XFILLER_0_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09476_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[13\]
+ net271 net291 net222 vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a211o_1
XANTENNA__06575__A _00754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06688_ _01223_ _01413_ _02324_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09492__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08427_ _03657_ _03755_ _03900_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__or3b_1
XFILLER_0_65_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05639_ _01350_ _01351_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08358_ net485 net416 _03719_ _03833_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload2 clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload2/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_22_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07309_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08289_ _03632_ _03661_ _03765_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ clknet_leaf_47_wb_clk_i net752 net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10251_ clknet_leaf_76_wb_clk_i _00243_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_104_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05638__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ clknet_leaf_9_wb_clk_i _00192_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05925__Y _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout250 _04729_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_2
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_4
Xfanout283 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\] vssd1
+ vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_4
Xfanout294 _03033_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07572__C net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10887__563 vssd1 vssd1 vccd1 vccd1 _10887__563/HI net563 sky130_fd_sc_hd__conb_1
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07494__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06049__A2 _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10518_ clknet_leaf_16_wb_clk_i _00386_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08205__A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10449_ clknet_leaf_47_wb_clk_i _00333_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05548__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05990_ net214 net184 _01663_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__a21oi_4
X_04941_ net441 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07660_ net131 _01676_ net167 _02835_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_49_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06611_ _02013_ _02073_ _02276_ _02282_ net254 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a221oi_4
X_07591_ net173 net144 _01658_ _03077_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__o31ai_1
X_09330_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ net6 _04312_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__a21oi_1
X_06542_ net119 net276 net111 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_66_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06395__A _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04908__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09261_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ _04459_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06473_ _02143_ _02145_ _02146_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__or3_1
XFILLER_0_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08212_ net462 _03689_ _03690_ _01283_ _03681_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__o32a_1
X_05424_ _01030_ _01048_ _01056_ _01034_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__a2bb2o_1
X_09192_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ _04407_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08143_ _00702_ _03628_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__or2_4
XFILLER_0_71_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05355_ net299 _01067_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout121_A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08074_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ net396 net298 net1004 _03589_ vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05286_ _00976_ _00997_ vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07025_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] net301 _00943_ _02679_
+ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout490_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] net797
+ net447 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__mux2_1
X_10914__659 vssd1 vssd1 vccd1 vccd1 net659 _10914__659/LO sky130_fd_sc_hd__conb_1
Xhold25 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05474__A team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold47 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__A2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold58 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ net299 _01665_ _03310_ _03481_ _03303_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__o32a_1
Xhold69 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06289__B net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07858_ net281 _03292_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__nand2_1
XANTENNA__07173__B1 _02673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06809_ _02479_ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__inv_2
X_07789_ _01050_ _01590_ _01598_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10661__RESET_B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09528_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] _00666_
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\] vssd1 vssd1
+ vccd1 vccd1 _04643_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09459_ net931 net208 _04601_ _04602_ vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__o22a_1
XFILLER_0_81_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07228__B2 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08025__A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10303_ clknet_leaf_47_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[16\]
+ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10234_ clknet_leaf_82_wb_clk_i net697 net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_10165_ clknet_leaf_7_wb_clk_i _00175_ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_10096_ clknet_leaf_80_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[1\]
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.labelPixel\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07164__B1 _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10998_ net392 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_44_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07467__A1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05478__B1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07758__B net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05140_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00853_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold506 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] vssd1 vssd1
+ vccd1 vccd1 net1176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05071_ _00672_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\] vssd1 vssd1
+ vccd1 vccd1 _00799_ sky130_fd_sc_hd__nor2_1
XANTENNA__09916__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_41_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08830_ _04173_ _04174_ net196 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07942__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08761_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ net235 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__mux2_1
X_05973_ net185 net176 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__nor2_2
X_07712_ _03260_ _03264_ _03267_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04924_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08692_ _01243_ _01251_ _04035_ _01250_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07643_ _01730_ _02765_ _03073_ _03105_ _03200_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__o32a_1
X_10983__624 vssd1 vssd1 vccd1 vccd1 _10983__624/HI net624 sky130_fd_sc_hd__conb_1
XFILLER_0_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06902__B1 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04909__Y _00651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07574_ _02033_ _02040_ net164 _02836_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_24_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09447__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09313_ net229 _04496_ _04497_ net405 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__a32o_1
XFILLER_0_119_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06525_ _02139_ _02195_ _02196_ _02198_ _02193_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__a311o_1
XFILLER_0_119_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout336_A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09244_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ _04444_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06456_ _02059_ _02072_ _02093_ _02128_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__o31a_1
XFILLER_0_17_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05407_ _01106_ _01107_ _01115_ _01060_ _01118_ vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09175_ net211 _04395_ _04397_ net402 net993 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__a32o_1
XFILLER_0_133_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06387_ net216 net175 net137 _01684_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__a31o_2
XANTENNA_fanout124_X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08126_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[9\]
+ _03612_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__or2_1
X_05338_ net397 _01049_ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ _03582_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ net297 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05269_ net427 _00979_ net426 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07008_ _02658_ _02667_ vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__xor2_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08959_ _04247_ net423 _04245_ vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10921_ net666 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XANTENNA__07697__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10852_ net528 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_67_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ clknet_leaf_66_wb_clk_i _00604_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08646__B1 _04070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07594__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10217_ clknet_leaf_0_wb_clk_i _00221_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10148_ clknet_leaf_1_wb_clk_i net751 net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10967__608 vssd1 vssd1 vccd1 vccd1 _10967__608/HI net608 sky130_fd_sc_hd__conb_1
X_10079_ clknet_leaf_28_wb_clk_i _00137_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_85_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07152__A3 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06310_ net441 net189 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07290_ _02921_ _02922_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[6\]
+ sky130_fd_sc_hd__or2_1
XANTENNA__06112__A1 _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06673__A _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06241_ _01672_ _01915_ _01917_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06392__B net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06172_ net215 net96 _01852_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold303 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[2\] vssd1
+ vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold314 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[5\] vssd1 vssd1 vccd1
+ vccd1 net984 sky130_fd_sc_hd__dlygate4sd3_1
X_05123_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] _00833_ vssd1 vssd1
+ vccd1 vccd1 _00836_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07612__A1 _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold325 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[1\] vssd1
+ vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 _00034_ vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold358 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ net892 net340 _01788_ _04905_ vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__a31o_1
Xhold369 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\] vssd1 vssd1
+ vccd1 vccd1 net1039 sky130_fd_sc_hd__dlygate4sd3_1
X_05054_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00780_ _00766_
+ vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09862_ _00726_ _03992_ _04804_ _04863_ _04861_ vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__a41o_1
XANTENNA__06179__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[11\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\]
+ _04160_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__or3_1
X_09793_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout286_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] net1074 net238 vssd1
+ vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__mux2_1
X_05956_ net134 net127 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_124_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04907_ net288 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _04075_ _04100_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__a21o_1
X_05887_ _00715_ _01575_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout453_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07626_ _02786_ _03169_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07557_ _01880_ _02743_ _03113_ _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06508_ net100 _02180_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07488_ net135 net142 _01729_ _01743_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09227_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ _04430_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__a21o_1
X_06439_ _01708_ _01732_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05199__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09158_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04379_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08109_ net943 _02672_ vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09089_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ _04328_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05927__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10002_ clknet_leaf_41_wb_clk_i _00022_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06477__B _01901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10904_ net570 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_15_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10835_ net511 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_137_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10766_ clknet_leaf_62_wb_clk_i _00587_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10697_ clknet_leaf_70_wb_clk_i _00528_ net350 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10251__Q team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05810_ _01494_ _01499_ _01500_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__o31a_2
X_06790_ _02410_ _02415_ _02460_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__and3_1
XANTENNA__05572__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05741_ _00774_ _00783_ _01442_ _00766_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[4\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06020__X _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08460_ _03753_ _03932_ _03927_ net130 vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__o211a_1
X_05672_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] _01260_
+ _01379_ _01380_ _01383_ vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__a2111o_1
X_07411_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] _02999_
+ net476 vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__o21ai_1
X_08391_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] _01259_ _01284_
+ _01305_ _03865_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__a41o_1
X_07342_ net476 net489 _00797_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07273_ _01389_ _02911_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[12\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_116_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ net251 _04275_ _04276_ net403 net874 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__a32o_1
X_06224_ net203 _01829_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__or2_2
XFILLER_0_54_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold100 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08389__A2 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06155_ net91 _01834_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout201_A _01517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold122 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05106_ net1006 _00817_ _00823_ net1065 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__a22o_1
Xhold144 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[8\] vssd1 vssd1
+ vccd1 vccd1 net814 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06086_ _01768_ _01769_ _01770_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__or3_1
Xhold155 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[14\]
+ vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[3\] vssd1 vssd1
+ vccd1 vccd1 net847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold188 team_07_WB.instance_to_wrap.ssdec_sdi vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__dlygate4sd3_1
X_05037_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__and4bb_1
X_09914_ net854 net154 net152 _04896_ vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold199 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[24\]
+ vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10434__RESET_B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07962__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input6_A gpio_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _04850_ _04851_ net1083 _04824_ vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_77_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10989__630 vssd1 vssd1 vccd1 vccd1 _10989__630/HI net630 sky130_fd_sc_hd__conb_1
XFILLER_0_119_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07681__B _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_77_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06988_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] _02651_
+ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__nand2_1
XANTENNA__06572__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06578__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ net1019 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net234 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05939_ _01628_ _01632_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08658_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04046_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07609_ _02254_ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__nor2_1
XANTENNA__05532__C1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08589_ _03606_ _04028_ net140 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__a21oi_1
X_10620_ clknet_leaf_48_wb_clk_i net870 net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06088__B1 _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10551_ clknet_leaf_20_wb_clk_i _00419_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10482_ clknet_leaf_22_wb_clk_i _00350_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06260__A0 _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09563__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10175__RESET_B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10104__RESET_B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__B1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06866__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10818_ net494 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10749_ clknet_leaf_68_wb_clk_i _00579_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10246__Q team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09568__A1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05838__Y _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07043__A2 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07960_ _01092_ net120 _03507_ _03508_ _03514_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_71_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06911_ _02497_ _02521_ _02578_ _02581_ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_71_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07891_ net259 _03316_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__or2_1
X_09630_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\] _04696_ net1075
+ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a21oi_1
X_06842_ net201 _02500_ _02512_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a21oi_1
X_09561_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ net795 net236 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__mux2_1
X_06773_ net428 net159 _01720_ _00672_ _01736_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__o221a_1
X_05724_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[20\]
+ _00824_ _00825_ net1011 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__a22o_1
X_08512_ _01793_ _03974_ _03966_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__o21ai_2
X_09492_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[18\]
+ net272 _04614_ _04621_ net221 vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__a221o_1
XANTENNA__07503__B1 _03050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08700__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05655_ _01364_ _01367_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__nor2_1
X_08443_ _03738_ _03916_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08374_ net488 _03849_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__nor2_1
XANTENNA__08059__B2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05586_ _01292_ _01294_ _01296_ _01298_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07325_ _02940_ _00974_ _00964_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout416_A team_07_WB.instance_to_wrap.team_07.heartPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07256_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06207_ _01887_ _01847_ _01827_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[0\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_115_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07187_ _02065_ net81 _02736_ _02831_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout204_X net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06138_ _01810_ _01814_ _01816_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10615__RESET_B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06069_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__or2_1
XANTENNA__08073__A_N net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout410 net412 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_2
Xfanout421 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] vssd1
+ vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout432 net433 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_2
Xfanout443 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[2\] vssd1 vssd1 vccd1
+ vccd1 net443 sky130_fd_sc_hd__clkbuf_2
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_1
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_4
Xfanout476 net484 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09828_ net971 _04836_ _04839_ _04824_ vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__o22a_1
Xfanout487 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__06545__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ net249 _04786_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05940__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10603_ clknet_leaf_47_wb_clk_i net910 net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout83 _02375_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_2
XFILLER_0_135_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout94 _01605_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_4
XFILLER_0_36_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09558__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07867__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10534_ clknet_leaf_21_wb_clk_i _00402_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06481__B1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10465_ clknet_leaf_14_wb_clk_i net729 net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_down
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06490__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10356__RESET_B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10396_ clknet_leaf_10_wb_clk_i net695 net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_92_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09722__A1 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ net642 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_126_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output45_A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06946__A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07113__Y _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05440_ _00964_ _01152_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05371_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] _00668_ _01067_
+ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_126_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07110_ _02033_ _02069_ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__or2_2
XFILLER_0_70_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05849__X _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08090_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[9\]
+ _00814_ net483 vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload20 clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_4
X_07041_ net156 _01700_ _01828_ net202 vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a31o_1
Xclkload31 clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_28_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload42 clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload53 clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__clkinv_8
Xclkload64 clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__inv_8
XANTENNA__10097__RESET_B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05297__A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload75 clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload86 clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__clkinv_8
X_08992_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_110_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07972__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10832__508 vssd1 vssd1 vccd1 vccd1 _10832__508/HI net508 sky130_fd_sc_hd__conb_1
X_07943_ _01068_ net162 _03309_ _03497_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__o211ai_1
XANTENNA__06399__Y _02073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout199_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10951__592 vssd1 vssd1 vccd1 vccd1 _10951__592/HI net592 sky130_fd_sc_hd__conb_1
X_07874_ _01051_ net118 net112 _01077_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09613_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\] _04664_ _04684_
+ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__or3_1
X_06825_ net433 net145 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout366_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09544_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[41\]
+ net225 _04605_ net879 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__a22o_1
X_06756_ net257 _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05707_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__nor2_1
X_06687_ _02354_ _02358_ _02359_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__or3b_1
X_09475_ net955 net207 _04610_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06575__B _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08426_ _03661_ net472 net468 vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__mux2_1
X_05638_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] vssd1 vssd1 vccd1
+ vccd1 _01351_ sky130_fd_sc_hd__and3b_1
XFILLER_0_18_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08357_ team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel team_07_WB.instance_to_wrap.team_07.flagPixel
+ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__or2_1
XANTENNA__08437__D1 _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05569_ net420 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 _01282_ sky130_fd_sc_hd__or3b_2
XFILLER_0_117_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload3 clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07308_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ _02930_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08288_ _00717_ net472 vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__nand2_1
XANTENNA__06591__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06463__B1 _02135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07239_ net129 net141 _02877_ _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__a31o_1
XANTENNA__10291__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10250_ clknet_leaf_82_wb_clk_i _00242_ net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05638__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10181_ clknet_leaf_8_wb_clk_i _00191_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05905__A_N _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06766__A1 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05935__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout240 net244 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_4
Xfanout251 _04270_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_2
Xfanout262 _01488_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_4
Xfanout273 _04591_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_4
Xfanout284 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\] vssd1
+ vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_4
Xfanout295 _03033_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07191__B2 _02842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07494__A2 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10517_ clknet_leaf_17_wb_clk_i _00385_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05829__B _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10448_ clknet_leaf_47_wb_clk_i _00332_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_110_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06006__A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05548__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10379_ clknet_leaf_15_wb_clk_i net694 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08221__A team_07_WB.instance_to_wrap.team_07.heartPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_04940_ net444 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
XANTENNA__06012__Y _01705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__B1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05980__A2 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05717__C1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07182__A1 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06610_ net254 _02275_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__or2_1
X_07590_ net87 _02109_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__nand2_1
XANTENNA__06676__A _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05580__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06541_ _01616_ _02213_ _02214_ _01618_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06395__B _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09260_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ net406 net230 _04460_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__a22o_1
X_06472_ _02139_ _02141_ _02078_ _02095_ _02118_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_138_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08211_ _01285_ _03684_ _03688_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__nor3_1
X_05423_ _01131_ _01133_ _01135_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__or3_1
X_09191_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ _04407_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08142_ _00702_ _03628_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__nor2_1
X_05354_ _00966_ _01048_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__or2_4
XANTENNA__08434__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08073_ net456 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__and2b_1
XFILLER_0_113_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05285_ _00976_ _00997_ vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout114_A _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07024_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\]
+ net449 vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08975_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\] net833
+ net447 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__mux2_1
Xhold15 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[0\]
+ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07018__Y _02673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07926_ _01084_ _01652_ _01700_ _03325_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__o211ai_1
Xhold48 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ _03410_ _03411_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06808_ net282 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1 vssd1
+ vccd1 vccd1 _02479_ sky130_fd_sc_hd__nand2_1
XANTENNA__06586__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07788_ _01590_ _01598_ _01050_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09527_ net921 net206 _04642_ vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06739_ net430 net431 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09458_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[4\]
+ net272 net220 vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09870__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08409_ _03810_ _03883_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ _01415_ _04549_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10630__RESET_B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07228__A2 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08025__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10302_ clknet_leaf_47_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[15\]
+ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08740__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06451__A3 _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ clknet_leaf_82_wb_clk_i net693 net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[3\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05936__Y _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10854__530 vssd1 vssd1 vccd1 vccd1 _10854__530/HI net530 sky130_fd_sc_hd__conb_1
X_10164_ clknet_leaf_8_wb_clk_i _00174_ net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05384__B _01005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10095_ clknet_leaf_82_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[0\]
+ net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.labelPixel\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07164__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05175__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10997_ net392 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_44_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07120__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold507 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\] vssd1 vssd1
+ vccd1 vccd1 net1177 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06007__Y _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05070_ net264 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ sky130_fd_sc_hd__inv_2
XFILLER_0_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05650__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08760_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] net1183 net237 vssd1
+ vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__mux2_1
X_05972_ net260 net176 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_81_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07711_ _02194_ _02219_ _02738_ _03044_ _03266_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__o221a_1
X_04923_ net2 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08691_ _01749_ _01755_ _04059_ _04111_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__or4_1
XANTENNA__07155__A1 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_10_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07642_ _01737_ _02261_ _03197_ _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07573_ net137 _01688_ net169 _03131_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_24_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09312_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04494_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06524_ net265 net87 _01711_ _02047_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__and4_1
XFILLER_0_119_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10429__Q team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_cleared vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ _04444_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06455_ net268 _02030_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__or2_2
XFILLER_0_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout329_A net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05406_ _01071_ _01103_ _01104_ _01075_ _01076_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__o32a_1
X_09174_ _04396_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06386_ _01680_ net166 _02057_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07030__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[8\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[7\] _03611_
+ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08958__A2 _01413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05337_ _00967_ _01048_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout117_X net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08056_ net455 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ net393 _03581_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05268_ net426 net428 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10838__514 vssd1 vssd1 vccd1 vccd1 _10838__514/HI net514 sky130_fd_sc_hd__conb_1
X_07007_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\]
+ _02649_ _02667_ _02668_ vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
X_05199_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] _00904_ vssd1 vssd1
+ vccd1 vccd1 _00912_ sky130_fd_sc_hd__xor2_1
XANTENNA__08591__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08958_ _01223_ _01413_ _00017_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__a21o_1
XANTENNA__07501__A_N net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08851__B1_N net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07909_ net259 _03370_ _03463_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__or3_1
X_08889_ _00708_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[1\]
+ net482 vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__o21a_1
XANTENNA__06587__Y _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ net665 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XANTENNA__05932__B _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07697__A2 _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851_ net527 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
X_10782_ clknet_leaf_66_wb_clk_i _00603_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06657__B1 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06409__B1 _02082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05379__B _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05947__X _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10895__652 vssd1 vssd1 vccd1 vccd1 net652 _10895__652/LO sky130_fd_sc_hd__conb_1
XFILLER_0_105_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05395__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10216_ clknet_leaf_86_wb_clk_i _00220_ net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ clknet_leaf_1_wb_clk_i net728 net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_89_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10078_ clknet_leaf_28_wb_clk_i _00136_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_85_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10249__Q team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06112__A2 _01789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__C_N net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06240_ _01851_ _01869_ _01902_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__and3b_1
XFILLER_0_127_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07121__Y _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06392__C _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06171_ net199 net92 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05122_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__or2_1
Xhold304 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[3\]
+ vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold315 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[8\] vssd1 vssd1
+ vccd1 vccd1 net985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold326 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold337 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_down vssd1
+ vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[7\] vssd1
+ vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09930_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\] _01786_
+ net155 net1025 vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__o31a_1
X_05053_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00763_ vssd1 vssd1
+ vccd1 vccd1 _00784_ sky130_fd_sc_hd__nand2_1
XANTENNA__06281__D1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold359 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\] vssd1 vssd1
+ vccd1 vccd1 net1029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09861_ _00762_ _04712_ _04862_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__or3b_1
XANTENNA__06179__A2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08812_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\] _04160_
+ net940 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__o21ai_1
X_09792_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[17\]
+ net238 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__mux2_1
X_05955_ net157 net149 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__nand2_4
XANTENNA__07128__A1 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07128__B2 _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A _00651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_04906_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] vssd1
+ vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _04053_ _04084_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_124_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05886_ _00715_ _01575_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__and2_1
X_07625_ net142 _03079_ _03182_ _03077_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__o22a_1
XANTENNA__10938__X net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07556_ _02235_ _03108_ _03109_ _01703_ _03112_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06507_ net100 _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__nor2_1
X_07487_ net184 _01744_ _02151_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09226_ _04435_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06438_ _02088_ _02110_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09157_ _04384_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06369_ _02037_ _02041_ _02034_ _02035_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08108_ _02672_ _03605_ vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08143__X _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09088_ _04333_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08039_ _03572_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ net394 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__mux2_1
XANTENNA__05927__B net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10001_ clknet_leaf_41_wb_clk_i _00021_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05007__X net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10903_ net569 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10834_ net510 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XANTENNA__05026__A_N net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07222__X _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10765_ clknet_leaf_66_wb_clk_i _00586_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10696_ clknet_leaf_70_wb_clk_i _00527_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05396__Y _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06014__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05369__B1 _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10733__RESET_B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05740_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] _00773_ vssd1
+ vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__or2_1
XANTENNA__05572__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05671_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\]
+ net420 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__or3b_1
XANTENNA__07530__A1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07410_ _02999_ _03000_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08390_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\] _03864_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07341_ _02945_ _02950_ _02952_ _02936_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[2\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07272_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ _02910_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09011_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__a31o_1
X_06223_ net202 _01829_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__nor2_2
XFILLER_0_60_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06154_ net91 _01834_ _01832_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold101 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[6\] vssd1
+ vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__A1 _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold123 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__dlygate4sd3_1
X_05105_ net481 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ _00821_ _00817_ net986 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__a32o_1
XFILLER_0_41_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__dlygate4sd3_1
X_06085_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] vssd1 vssd1 vccd1 vccd1
+ _01770_ sky130_fd_sc_hd__or3b_1
XFILLER_0_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold145 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[2\] vssd1 vssd1
+ vccd1 vccd1 net837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05036_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[5\]
+ _00767_ vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__nor3_1
X_09913_ _01781_ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__nand2_1
Xhold178 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[12\] vssd1 vssd1
+ vccd1 vccd1 net848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[2\]
+ vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout396_A _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09844_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\] _04848_ net269
+ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07962__B _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09775_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__or4bb_1
XANTENNA__07681__C _03144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06987_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] _02650_
+ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__and2_1
XANTENNA__06578__B net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout184_X net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08726_ net885 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05938_ _00754_ _01631_ net100 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_1_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08657_ _00707_ _04050_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05869_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] net178
+ _01547_ net158 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07608_ _01811_ net165 _01672_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08588_ net801 net730 vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__nand2_1
XANTENNA__06594__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07042__X _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07539_ _02080_ _02129_ _02150_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__a21o_2
XFILLER_0_9_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10550_ clknet_leaf_19_wb_clk_i _00418_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09209_ _04420_ _04422_ _04421_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10481_ clknet_leaf_22_wb_clk_i _00349_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06260__A1 _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout97_X net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07760__A1 _01067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05392__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__B2 _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05960__X _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10817_ net493 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08068__A2 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10748_ clknet_leaf_68_wb_clk_i _00578_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08473__C1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06009__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10679_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[11\]
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08224__A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06787__C1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06910_ _02579_ _02580_ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07890_ _03442_ _03443_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__nand2_1
XANTENNA__06003__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05583__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06841_ net217 _02511_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__nor2_1
XANTENNA__06031__X _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09560_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ net809 net236 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__mux2_1
X_06772_ net93 _02414_ _02416_ net108 _02443_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__a221o_1
X_08511_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__inv_2
X_05723_ net989 _00824_ _00825_ net1102 _01430_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__a221o_1
X_09491_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _04613_ _04616_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__nand3_1
XANTENNA__07503__A1 _03058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08442_ net459 _03915_ _03695_ _03694_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__o211a_1
X_05654_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] _01301_
+ _01362_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08373_ team_07_WB.instance_to_wrap.team_07.buttonPixel _03700_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05585_ _01286_ _01289_ _01291_ _01281_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout144_A _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07324_ _02939_ _00973_ _01109_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10437__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07255_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout311_A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06206_ _01851_ _01869_ _01876_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__or4_1
X_07186_ _02835_ _02837_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06137_ net289 net132 net127 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__a211o_1
XANTENNA__10814__D team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11017__642 vssd1 vssd1 vccd1 vccd1 _11017__642/HI net642 sky130_fd_sc_hd__conb_1
XFILLER_0_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06068_ _01750_ _01751_ _01753_ _01754_ _01752_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout400 net410 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_2
Xfanout411 net412 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout422 net423 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_2
XFILLER_0_10_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05019_ net280 _00752_ vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__nor2_2
Xfanout433 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\] vssd1 vssd1 vccd1
+ vccd1 net433 sky130_fd_sc_hd__buf_2
XANTENNA__06589__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout444 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\] vssd1 vssd1 vccd1
+ vccd1 net444 sky130_fd_sc_hd__buf_2
Xfanout455 net456 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_2
Xfanout466 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.frameBufferLowNibble
+ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_4
Xfanout477 net484 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_2
X_09827_ _00657_ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__nor2_1
Xfanout488 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_2
XANTENNA__06545__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ _04767_ _04786_ _04787_ net249 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08709_ _04126_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ _04115_ vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__mux2_1
X_09689_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\]
+ _04736_ _00655_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05940__B net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07213__A _02073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10602_ clknet_leaf_47_wb_clk_i net894 net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout84 _02177_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout95 net97 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10533_ clknet_leaf_21_wb_clk_i _00401_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05939__Y _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06481__A1 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ clknet_leaf_13_wb_clk_i net742 net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_up
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05387__B _01014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10395_ clknet_leaf_10_wb_clk_i _00039_ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06233__B2 _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11016_ net391 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08930__A0 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08446__C1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05370_ net437 _00668_ _01067_ vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__o21a_2
XFILLER_0_43_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload10 clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_12
Xclkload21 clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_12
X_07040_ _02214_ _02258_ _02692_ _02694_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload32 clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__inv_6
XANTENNA__08749__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload43 clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__inv_16
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload54 clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload65 clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__inv_8
Xclkload76 clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_73_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload87 clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__inv_8
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07793__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__and4_1
XFILLER_0_76_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07972__A1 _01113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07942_ _01068_ net161 _01653_ _01083_ _01699_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__a221o_1
X_10871__547 vssd1 vssd1 vccd1 vccd1 _10871__547/HI net547 sky130_fd_sc_hd__conb_1
X_07873_ _01051_ net118 _03427_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__o21a_1
X_09612_ _04664_ _04684_ net1052 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__o21ai_1
X_06824_ net433 net145 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09543_ net879 net224 _04605_ net916 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06755_ _00671_ _00985_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout261_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout359_A net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05706_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__or2_1
X_09474_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[12\]
+ net271 net291 net222 vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a211o_1
X_06686_ _02338_ _02345_ _02346_ _02355_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__and4_1
X_08425_ _03638_ _03641_ net467 vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__or3b_1
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05637_ net421 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] vssd1 vssd1 vccd1
+ vccd1 _01350_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08356_ _03828_ _03829_ _03831_ _03629_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06872__A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05568_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\]
+ _00677_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__or3_2
XFILLER_0_117_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload4 clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__10167__Q team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08988__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07307_ _02930_ _02933_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[0\]
+ sky130_fd_sc_hd__or2_1
X_08287_ net468 _03642_ _03639_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05499_ net422 _00692_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__or3_1
XANTENNA__06591__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05266__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07238_ net121 _01936_ _02861_ _02873_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__nor4_1
XFILLER_0_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07169_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] net301 net300 team_07_WB.instance_to_wrap.team_07.label_num_bus\[28\]
+ _02820_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10180_ clknet_leaf_8_wb_clk_i _00190_ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05935__B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout230 _04427_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__buf_2
Xfanout241 net242 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
Xfanout252 _04270_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_2
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_4
Xfanout274 _01622_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07715__A1 _00754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout285 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\] vssd1
+ vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_2
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07191__A2 _02838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05951__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09142__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07494__A3 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05398__A _01000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10516_ clknet_leaf_17_wb_clk_i _00384_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10447_ clknet_leaf_54_wb_clk_i _00331_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06006__B net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10378_ clknet_leaf_15_wb_clk_i _00037_ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_23_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07954__A1 _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06022__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__A1 _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10147__SET_B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07182__A2 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10309__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06390__B1 _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06676__B _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06540_ net267 net276 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_66_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06471_ _02064_ _02144_ _02137_ _02142_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__or4b_1
XFILLER_0_75_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08063__A_N net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08210_ _03688_ _03685_ _03687_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__and3b_1
X_05422_ _01007_ _01134_ _01107_ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__or3b_1
X_09190_ net211 _04406_ _04408_ net404 net1028 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08141_ net54 net52 vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05353_ _00966_ _01048_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08434__A2 _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08072_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ _03576_ net456 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05284_ net429 net430 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07023_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] _00829_ _00942_
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\] vssd1 vssd1 vccd1 vccd1
+ _02678_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08974_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] net825
+ net447 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__mux2_1
Xhold16 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold27 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07028__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07925_ _03320_ _03476_ _03478_ _03479_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__a211o_1
Xhold38 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07856_ _01678_ _03321_ _03326_ _01689_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06867__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06807_ _02468_ _02469_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__or2_1
X_07787_ _01056_ _01597_ _01604_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__and3_1
X_04999_ net39 net38 net10 net9 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__or4_1
XANTENNA__06586__B _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[32\]
+ net270 _04641_ net291 net223 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__a221o_1
X_06738_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ net430 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09457_ net417 _01416_ _04589_ net290 vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__o31a_1
X_06669_ _02340_ _02341_ _02339_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06133__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09870__A1 _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ _03808_ _03882_ net487 vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09388_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\] vssd1
+ vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08339_ net474 _03639_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10301_ clknet_leaf_47_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[14\]
+ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10670__RESET_B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10958__599 vssd1 vssd1 vccd1 vccd1 _10958__599/HI net599 sky130_fd_sc_hd__conb_1
X_10232_ clknet_leaf_82_wb_clk_i net714 net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[2\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10163_ clknet_leaf_8_wb_clk_i _00173_ net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input37_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ clknet_leaf_33_wb_clk_i team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[3\]
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05952__Y _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06496__B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10996_ net392 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07120__B _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07624__B1 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06017__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold508 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\] vssd1 vssd1
+ vccd1 vccd1 net1178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07927__A1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07119__Y _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05971_ net178 net158 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__nor2_4
X_07710_ _01729_ _02277_ _03206_ _03265_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__a211o_1
X_04922_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
X_08690_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01757_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07641_ _01722_ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__nand2_1
XANTENNA__06902__A2 _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07572_ net137 net105 net167 vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_105_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_50_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09311_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[11\]
+ _04494_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06523_ net98 net93 _02176_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__or3b_1
XFILLER_0_8_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09242_ net231 _04446_ _04447_ net407 net1084 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__a32o_1
XFILLER_0_119_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06454_ net268 _02030_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__nor2_2
XANTENNA__06666__B2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04935__A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05405_ _00669_ _01020_ _01061_ _01069_ vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__o22a_1
X_09173_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04391_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__and3_1
X_06385_ net129 _01676_ net166 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08124_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[6\]
+ _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06418__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07030__B _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05336_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] _00669_ vssd1
+ vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__nand2_2
X_10920__665 vssd1 vssd1 vccd1 vccd1 net665 _10920__665/LO sky130_fd_sc_hd__conb_1
XFILLER_0_126_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08055_ net456 net452 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__and3b_1
X_05267_ net426 _00671_ _00979_ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10877__553 vssd1 vssd1 vccd1 vccd1 _10877__553/HI net553 sky130_fd_sc_hd__conb_1
X_07006_ _02651_ _02659_ _02664_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05198_ _00909_ _00910_ _00908_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__a21o_1
XANTENNA__07918__A1 _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10010__RESET_B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05916__D net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08957_ _04246_ net425 _04245_ vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__mux2_1
X_07908_ _03369_ _03462_ _03368_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__a21oi_1
X_08888_ _00708_ _01429_ _04209_ net1086 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__a22o_1
XANTENNA__06597__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07839_ _03393_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__inv_2
XANTENNA__06354__B1 _02027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ net526 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XANTENNA__06519__A1_N _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09509_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[25\]
+ net271 _04584_ net224 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__a211o_1
X_10781_ clknet_leaf_66_wb_clk_i _00602_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07221__A _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06409__B2 _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07082__A1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10215_ clknet_leaf_0_wb_clk_i _00219_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09435__X _04584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07891__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ clknet_leaf_1_wb_clk_i net780 net308 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10077_ clknet_leaf_28_wb_clk_i _00135_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06300__A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06345__B1 _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload2_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06794__X team_07_WB.instance_to_wrap.team_07.recPLAYER.playerDetect vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10979_ net620 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_84_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06648__A1 _02080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06648__B2 _02135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07131__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06170_ _01839_ _01842_ _01850_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__and3b_1
XFILLER_0_108_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05121_ _00833_ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold305 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[16\]
+ vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold327 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[13\] vssd1 vssd1
+ vccd1 vccd1 net997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold349 team_07_WB.instance_to_wrap.team_07.label_num_bus\[1\] vssd1 vssd1 vccd1
+ vccd1 net1019 sky130_fd_sc_hd__dlygate4sd3_1
X_05052_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00655_ _00761_
+ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__and3_1
XANTENNA__06820__A1 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06820__B2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09860_ _00652_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _00772_
+ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__or3_1
XFILLER_0_110_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08811_ _04161_ _04162_ net195 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__a21oi_1
X_09791_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] _04808_ _04811_
+ _04813_ vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__a22o_1
X_08742_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[16\]
+ net238 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05954_ net160 net145 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08673_ _04080_ _04098_ _04084_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_124_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06210__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05885_ _01574_ _01575_ _00715_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout174_A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07624_ _01666_ _01734_ _02278_ _03120_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_36_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07555_ _01666_ _03077_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout341_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06506_ net284 net92 _01609_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07486_ _01715_ _02045_ _03046_ _01714_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__and4b_1
XFILLER_0_9_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09225_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ _04430_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__and3_1
X_06437_ _02110_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09156_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04379_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06368_ net170 _02040_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__nand2_1
XANTENNA__06880__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09053__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08107_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] _02671_
+ net1087 vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05319_ _01029_ _01020_ _01024_ _01031_ vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__and4b_1
X_09087_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ _04328_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__and3_1
X_06299_ _01401_ net441 net438 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08038_ _00706_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ net396 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06811__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10000_ clknet_leaf_41_wb_clk_i net1046 net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout87_A _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ clknet_leaf_42_wb_clk_i _00029_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09513__B1 _04584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10902_ net568 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_0_98_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10833_ net509 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_15_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10764_ clknet_leaf_66_wb_clk_i _00585_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10695_ clknet_leaf_70_wb_clk_i _00526_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07886__A _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10973__614 vssd1 vssd1 vccd1 vccd1 _10973__614/HI net614 sky130_fd_sc_hd__conb_1
XFILLER_0_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06566__B1 _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ clknet_leaf_36_wb_clk_i _00167_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06581__A3 _02254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06030__A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08858__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05670_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\]
+ net420 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_102_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07530__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07340_ _01175_ _02417_ _02951_ _00965_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07271_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__a21oi_1
X_09010_ _04274_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__inv_2
X_06222_ net156 _01736_ _01828_ net202 vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a31o_2
XANTENNA__07796__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07046__A1 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06153_ net103 _01828_ _01833_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold102 _00111_ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08404__B _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05104_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[13\]
+ _00824_ _00825_ net1016 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__a22o_1
Xhold124 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[3\] vssd1 vssd1
+ vccd1 vccd1 net794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__dlygate4sd3_1
X_06084_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold146 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold157 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[12\]
+ vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\] vssd1 vssd1
+ vccd1 vccd1 net838 sky130_fd_sc_hd__dlygate4sd3_1
X_05035_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__or4bb_1
X_09912_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[15\] _01780_
+ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__nand2_1
Xhold179 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[5\] vssd1 vssd1
+ vccd1 vccd1 net849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09843_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\]
+ _04844_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__and3_1
XANTENNA__06557__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09774_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__or4_1
X_06986_ _00713_ _02648_ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__nor2_1
XANTENNA__06578__C net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05937_ net94 net86 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__nand2_1
X_08725_ _04134_ _04137_ _04136_ vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_1_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08849__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout177_X net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ _01249_ _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__and2_1
X_05868_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] _01546_
+ _01561_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__and3_1
XANTENNA__06875__A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ net188 _02073_ _02744_ _02863_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__a211oi_2
X_08587_ net730 net140 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__nor2_1
XANTENNA__05532__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05799_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\]
+ _01486_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__nand3_1
XFILLER_0_37_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07538_ _03091_ _03096_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_944 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07469_ net413 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ _03024_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09208_ _04418_ _04419_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10480_ clknet_leaf_22_wb_clk_i _00348_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09139_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ _04370_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06115__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05954__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07760__A2 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10342__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06720__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05523__B2 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10816_ clknet_leaf_89_wb_clk_i _00036_ _00066_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10747_ clknet_leaf_68_wb_clk_i _00577_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06009__B net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05826__A2 _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10678_ clknet_leaf_59_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[10\]
+ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10823__499 vssd1 vssd1 vccd1 vccd1 _10823__499/HI net499 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_58_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06025__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06787__B1 _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07200__A1 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06003__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07127__Y _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ net432 _00694_ _02510_ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__o21a_1
XANTENNA__07200__B2 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06771_ net108 _02416_ _02441_ net116 _02442_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08510_ _03966_ _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__nand2_2
X_05722_ net483 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09490_ net904 net208 _04620_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08441_ net460 _03914_ _03676_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05653_ _01349_ _01364_ _01365_ _01347_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08372_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03847_ _00727_
+ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05584_ _01295_ _01296_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07323_ net427 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout137_A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07254_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ _02896_ _02899_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[6\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07019__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06205_ _01878_ _01885_ net96 vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07185_ _01732_ _02836_ _01725_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06136_ _01808_ _01810_ _01815_ _01816_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06778__B1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06067_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__nand2_1
Xfanout401 net410 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_2
Xfanout412 _00807_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_8
X_05018_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] net288
+ vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_6_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout423 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[1\] vssd1
+ vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06222__X _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout434 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[0\] vssd1 vssd1 vccd1
+ vccd1 net434 sky130_fd_sc_hd__buf_4
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout445 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[0\] vssd1 vssd1 vccd1
+ vccd1 net445 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06589__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout456 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_4
Xfanout467 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[3\] vssd1
+ vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_2
X_09826_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[6\] _04833_ vssd1 vssd1
+ vccd1 vccd1 _04838_ sky130_fd_sc_hd__and4_1
Xfanout478 net479 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_4
Xfanout489 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_2
XANTENNA__05202__B1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\] _04783_ vssd1
+ vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_5_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_06969_ _02562_ _02631_ _02636_ _02639_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_69_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08708_ net263 _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__and2_1
X_09688_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] _04738_ _04739_
+ _04734_ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09495__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08639_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_90_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05014__A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10601_ clknet_leaf_47_wb_clk_i _00465_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout85 _02177_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10532_ clknet_leaf_25_wb_clk_i _00400_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05949__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout96 net97 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_2
XFILLER_0_80_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10463_ clknet_leaf_22_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_select
+ net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06481__A2 _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05020__Y _00754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ clknet_leaf_11_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[2\]
+ net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05955__Y _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11015_ net641 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XANTENNA__09443__X _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08446__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10979__620 vssd1 vssd1 vccd1 vccd1 _10979__620/HI net620 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_136_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload11 clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinv_8
Xclkload22 clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_12
Xclkload33 clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__clkinv_4
Xclkbuf_leaf_75_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xclkload44 clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__inv_8
Xclkload55 clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__inv_8
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload66 clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload66/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload77 clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_73_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload88 clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07793__B _01069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ _04258_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_110_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07972__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07941_ net259 _03310_ _03324_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__nor3_1
X_07872_ net286 _01115_ _03390_ _03394_ _03288_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__a311o_1
XANTENNA__05881__X _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ _04666_ _04683_ _04684_ _04664_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__a32o_1
X_06823_ net95 _02471_ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09542_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[39\]
+ net224 _04605_ net839 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__a22o_1
X_06754_ net217 _02418_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05705_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07488__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06685_ _02079_ net84 _02329_ _02357_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__a31o_1
X_09473_ net934 net207 _04609_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout254_A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ net475 _03640_ net469 vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a21oi_2
X_05636_ _01348_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10448__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08355_ net472 _03631_ _03659_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05567_ _01278_ _01279_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__nor2_1
XANTENNA__04944__Y _00684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07306_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ _02932_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__a21oi_1
Xclkload5 clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_8
X_08286_ _03763_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05498_ net422 _00692_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07237_ _01743_ _02758_ _02887_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__and3_1
XANTENNA__07660__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07168_ net450 team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\] net398 vssd1
+ vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06119_ _01723_ _01797_ _01799_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a21bo_1
X_07099_ _02739_ _02751_ _02752_ _02748_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout220 net221 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
Xfanout231 _04427_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_2
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout253 _02170_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
Xfanout264 _00798_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_4
XANTENNA__07176__B1 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 _01622_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_2
XANTENNA__07715__A2 _01961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout286 net287 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_4
Xfanout297 _03026_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_2
X_09809_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\] net269 _04826_
+ vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__o21ba_1
XANTENNA__05951__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09468__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08676__B1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05015__Y _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10515_ clknet_leaf_18_wb_clk_i _00383_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07651__A1 _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10446_ clknet_leaf_39_wb_clk_i _00330_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10377_ clknet_leaf_11_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[2\]
+ net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07954__A2 _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06303__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07118__B _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07167__B1 _02673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__S net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07706__A2 _01901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08667__B1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06470_ net283 _01621_ _02104_ _02100_ net265 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a32o_1
XANTENNA__06142__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05421_ _01061_ _01079_ _01097_ _01103_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_138_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08419__B1 _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08140_ _02670_ net146 vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05589__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05352_ _00669_ _00967_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08071_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ _03575_ net456 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07642__A1 _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05283_ _00993_ _00995_ vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__nand2_1
X_07022_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] _00829_ _02676_
+ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_112_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08973_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] net819
+ net448 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__mux2_1
Xhold17 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold28 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07028__B _00754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07924_ _03313_ _03315_ net256 vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__o21ai_1
Xhold39 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ net274 _03294_ _03299_ _03300_ _03285_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__o32a_1
XFILLER_0_78_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06905__B1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06806_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] _02467_ _02476_
+ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a21bo_1
X_04998_ net19 net8 net33 net30 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__or4_1
X_07786_ _01597_ _01604_ _01056_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07044__A _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09525_ _01420_ _04640_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__or3b_1
X_06737_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ net430 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06668_ net99 _01616_ _02312_ _02332_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06133__A1 _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ net911 net208 _04600_ vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__o21a_1
XANTENNA__06883__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09870__A2 _01789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ _03707_ _03709_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__o21ai_1
X_05619_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ net445 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__mux2_1
X_06599_ net262 _01720_ _02271_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a21oi_1
X_09387_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ _01475_ _02984_ _04548_ vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__o22a_1
X_08338_ net470 net467 vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07633__A1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08269_ _03739_ _03747_ _03723_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08830__B1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10300_ clknet_leaf_47_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[13\]
+ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05011__B net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10231_ clknet_leaf_88_wb_clk_i net453 net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_30_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10162_ clknet_leaf_3_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[9\]
+ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10093_ clknet_leaf_58_wb_clk_i team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[2\]
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05962__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07164__A3 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10995_ net636 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_26_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07872__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10816__Q net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06017__B net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05696__X _01409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold509 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[0\] vssd1 vssd1
+ vccd1 vccd1 net1179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10429_ clknet_leaf_31_wb_clk_i _00313_ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_cleared
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10727__RESET_B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07927__A2 _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05938__A1 _00754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06033__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05970_ net261 _01657_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__nor2_4
XFILLER_0_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_04921_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05591__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07640_ _01645_ _02744_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__nor2_2
XFILLER_0_73_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07571_ _01680_ net167 _01739_ net170 vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09310_ net229 _04493_ _04495_ net404 net1132 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__a32o_1
X_06522_ net97 net89 _02176_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_24_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09241_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ _04444_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__nand2_1
X_06453_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] _02030_
+ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_90_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05404_ _01057_ _01059_ _01070_ _00967_ _01116_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__o221a_1
X_09172_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04391_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__a21o_1
X_06384_ _01675_ _02056_ _02054_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_69_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[5\]
+ _03609_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__or2_1
XANTENNA__06418__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05335_ _00668_ net436 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__nor2_4
XFILLER_0_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07030__C _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout217_A _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08054_ net1137 net296 _03580_ vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__a21o_1
X_05266_ net429 net430 _00978_ _00975_ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07005_ _02660_ _02664_ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05197_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00904_ vssd1 vssd1
+ vccd1 vccd1 _00910_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07918__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10461__Q team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08956_ net476 net425 vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_129_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05782__A _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07907_ _01057_ net178 vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08887_ _03591_ _03592_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__mux2_2
XANTENNA__06597__B _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ net277 _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__or2_1
X_07769_ _03316_ _03322_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09508_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[25\]
+ net222 _04605_ net869 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__a22o_1
X_10780_ clknet_leaf_65_wb_clk_i _00601_ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09439_ net220 _04587_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07221__B _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06118__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05022__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05957__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07082__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06405__X _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10214_ clknet_leaf_86_wb_clk_i _00218_ net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10145_ clknet_leaf_1_wb_clk_i net758 net308 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10076_ clknet_leaf_35_wb_clk_i _00134_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10599__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10978_ net619 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_58_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07131__B net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06028__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09598__A1 _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05120_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold306 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\] vssd1 vssd1
+ vccd1 vccd1 net976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold317 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\] vssd1 vssd1
+ vccd1 vccd1 net987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold328 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\] vssd1 vssd1
+ vccd1 vccd1 net998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 _00103_ vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__dlygate4sd3_1
X_05051_ _00781_ _00782_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\]
+ _00766_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[6\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_22_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08810_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\] _04160_
+ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__or2_1
X_09790_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] _04810_ vssd1
+ vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06584__A1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08741_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ net234 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__mux2_1
X_05953_ _01643_ _01645_ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_107_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08672_ _04092_ _04089_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__and2b_1
X_05884_ _01574_ _01575_ _00715_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_124_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07623_ _02067_ _02150_ _03149_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07554_ net141 _03077_ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__or2_1
XANTENNA__04946__A team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06505_ _02109_ _02163_ _02169_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10844__520 vssd1 vssd1 vccd1 vccd1 _10844__520/HI net520 sky130_fd_sc_hd__conb_1
X_07485_ _01903_ _02040_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout334_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09224_ net231 _04433_ _04434_ net408 net1128 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09038__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06436_ _01680_ net168 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__and2_2
XFILLER_0_17_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09155_ net210 _04382_ _04383_ net401 net1064 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06367_ net131 net124 net170 net141 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__and4_1
XANTENNA__10649__RESET_B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout122_X net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08106_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] _02671_
+ vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05318_ net194 _01014_ _01021_ _01030_ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__o31a_1
XFILLER_0_114_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06298_ net177 _01973_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__xnor2_1
X_09086_ net212 _04331_ _04332_ net399 net1080 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__a32o_1
XANTENNA__06272__B1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08037_ net456 net452 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__and3b_1
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05249_ _00957_ _00958_ _00961_ vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ clknet_leaf_42_wb_clk_i net1012 net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_08939_ net491 _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__nor2_1
XANTENNA__08316__A2 _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10931__581 vssd1 vssd1 vccd1 vccd1 _10931__581/HI net581 sky130_fd_sc_hd__conb_1
XFILLER_0_93_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10901_ net567 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_84_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10832_ net508 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_15_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07232__A _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10763_ clknet_leaf_62_wb_clk_i _00584_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10694_ clknet_leaf_70_wb_clk_i _00525_ net350 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05958__Y _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07886__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06566__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ clknet_leaf_36_wb_clk_i net802 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06311__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ clknet_leaf_30_wb_clk_i _00117_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06030__B _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_102_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10828__504 vssd1 vssd1 vccd1 vccd1 _10828__504/HI net504 sky130_fd_sc_hd__conb_1
XANTENNA__07530__A3 _02082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06029__Y _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07270_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06221_ net176 net157 vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__nand2_4
XANTENNA__10614__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06152_ _01644_ net102 net197 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07046__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold103 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[3\] vssd1
+ vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__dlygate4sd3_1
X_05103_ net482 _00814_ _00822_ vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__and3_2
Xhold114 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[4\] vssd1 vssd1
+ vccd1 vccd1 net784 sky130_fd_sc_hd__dlygate4sd3_1
X_06083_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__or2_1
Xhold125 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[6\] vssd1 vssd1
+ vccd1 vccd1 net806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold147 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[2\]
+ vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[1\] vssd1 vssd1
+ vccd1 vccd1 net828 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ net852 net154 net152 _04894_ vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__a22o_1
X_05034_ _00763_ _00765_ vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__nand2_2
Xhold169 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[38\]
+ vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_81_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10764__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09842_ net1078 _04847_ _04849_ net247 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__o22a_1
XFILLER_0_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06557__A1 _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\] _01769_ _04797_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] vssd1 vssd1 vccd1 vccd1
+ _04798_ sky130_fd_sc_hd__or4b_1
XANTENNA__06221__A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06985_ _02647_ _02648_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout284_A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08724_ _01240_ _04080_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__and2_1
X_05936_ net115 net108 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__nand2_2
XANTENNA__06309__A1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _04073_ _04082_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout451_A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05867_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] net162
+ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__xnor2_4
X_07606_ _03078_ _03164_ _03159_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.boomGen.boomDetect
+ sky130_fd_sc_hd__a21o_1
X_08586_ net146 _04027_ _03965_ vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05798_ _01490_ _01491_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_49_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07537_ net124 net144 _03079_ _03095_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__or4b_1
XFILLER_0_64_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07809__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07809__B2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07468_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ net294 _03035_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[29\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09207_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[16\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__o2111ai_2
XANTENNA__06493__B1 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06419_ _02074_ _02092_ _02090_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a21o_1
XANTENNA__05778__Y _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07399_ _02992_ _02993_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09138_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04369_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__o31a_1
XANTENNA__10412__RESET_B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09069_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ _04318_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__o31a_1
XFILLER_0_124_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05794__X _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05954__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06548__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06548__B2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06131__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05018__Y _00752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05970__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06720__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10815_ clknet_leaf_7_wb_clk_i team_07_WB.instance_to_wrap.team_07.recHEART.heartDetect
+ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.heartPixel sky130_fd_sc_hd__dfrtp_4
XFILLER_0_138_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10746_ clknet_leaf_67_wb_clk_i _00576_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06484__B1 _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10677_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[9\]
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05588__A_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06025__B net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07200__A2 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06041__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ _02417_ _02440_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__nand2_1
X_05721_ net481 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ _00822_ _00824_ net986 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__a32o_1
XFILLER_0_78_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07503__A3 _03062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08440_ _00731_ _03913_ _03679_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__a21oi_1
X_05652_ _01331_ _01337_ _01342_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__or3b_1
XFILLER_0_59_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06711__A1 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08371_ _03777_ _03779_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__a21oi_1
X_05583_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] vssd1 vssd1 vccd1
+ vccd1 _01296_ sky130_fd_sc_hd__or3b_2
XFILLER_0_129_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07322_ _00672_ _02938_ _02937_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07253_ _00718_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06204_ net94 _01879_ _01883_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07184_ _01715_ _01873_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__nor2_4
XFILLER_0_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_3_0_wb_clk_i_X clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06135_ net285 _01812_ _01813_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__nand3_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06066_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout402 net410 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_2
X_05017_ _00635_ _00649_ vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__nor2_1
XANTENNA__05450__B2 _01069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout413 _00706_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout424 net425 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_2
Xfanout435 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[2\] vssd1 vssd1
+ vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_4
Xfanout446 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[0\] vssd1 vssd1 vccd1
+ vccd1 net446 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input4_A gpio_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ net1047 _04834_ _04837_ vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__o21a_1
XANTENNA__07047__A _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_2
Xfanout468 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[3\] vssd1
+ vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout479 net480 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout287_X net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\] _04783_ vssd1
+ vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__nand2_1
X_06968_ _02556_ _02637_ _02638_ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__a21o_1
XANTENNA__06886__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ _01238_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__a41o_1
X_05919_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] _01593_
+ _01580_ _01578_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__o2bb2a_1
X_09687_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] _04738_ vssd1
+ vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06899_ net288 _02568_ _02562_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__o21ba_1
X_08638_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ net457 _04062_ _04063_ _04065_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__o311a_1
XFILLER_0_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08569_ _04015_ _04016_ _03996_ vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__o21a_1
XANTENNA__07213__C _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10600_ clknet_leaf_54_wb_clk_i _00464_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05014__B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout86 _01629_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_4
XFILLER_0_65_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10531_ clknet_leaf_25_wb_clk_i _00399_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout97 _01601_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__buf_2
XANTENNA__05949__B _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05301__Y _01014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10462_ clknet_leaf_13_wb_clk_i net1002 net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05668__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10393_ clknet_leaf_11_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[1\]
+ net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05965__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06413__X _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11014_ net390 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XANTENNA__05971__Y _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10729_ clknet_leaf_79_wb_clk_i _00559_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload12 clknet_leaf_88_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__inv_12
XANTENNA__06036__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload23 clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__clkinv_8
Xclkload34 clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__clkinv_2
Xclkload45 clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload56 clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_114_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload67 clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_24_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload78 clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_16
XTAP_TAPCELL_ROW_114_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07940_ _01067_ net219 _03314_ _03494_ net257 vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_110_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07709__B1 _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06042__Y _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_44_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07871_ _03421_ _03422_ _03340_ _03346_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__a211o_1
XANTENNA__07185__A1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\] _04682_ vssd1
+ vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__nand2_1
X_06822_ net95 _02471_ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__and2_1
X_09541_ _04651_ net839 net224 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__mux2_1
X_06753_ _00973_ net201 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05704_ net417 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ _01415_ vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__or3_1
XANTENNA__07488__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09472_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[11\]
+ net273 net293 net224 vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a211o_1
X_06684_ _02336_ _02349_ _02352_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__and3b_1
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09882__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08423_ net784 _03897_ _03653_ vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05635_ net420 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 _01348_ sky130_fd_sc_hd__and3b_1
XFILLER_0_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08354_ _03632_ _03637_ _03766_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_135_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05566_ _01270_ _01272_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07305_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_22_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08285_ net467 _03641_ _03660_ _03667_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__o311a_1
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05497_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ _01201_ _01208_ _01209_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__or4b_1
Xclkload6 clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA_fanout414_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07236_ net171 _02082_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07660__A2 _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07167_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] net302 _02673_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout202_X net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06118_ net199 _01798_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07098_ net144 _01669_ _01664_ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a21o_1
X_06049_ net176 _01737_ net185 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout210 _04376_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_2
Xfanout221 _04582_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout232 _03594_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_4
Xfanout243 net244 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_2
Xfanout254 net256 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07176__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_4
Xfanout276 _01620_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_4
X_09808_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\] _04825_ vssd1
+ vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__and2_1
Xfanout287 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\] vssd1
+ vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_4
Xfanout298 _03026_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06923__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\] _04772_ vssd1
+ vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05025__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08055__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10514_ clknet_leaf_18_wb_clk_i _00382_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08770__S net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07651__A2 _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05966__Y _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10445_ clknet_leaf_39_wb_clk_i _00329_ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07939__B1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05695__A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10376_ clknet_leaf_11_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[1\]
+ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06611__B1 _02276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05982__X _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09998__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05717__A2 _01413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07702__X _03258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09987__D net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05420_ _01026_ _01110_ _01132_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07150__A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05351_ net435 net397 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__nor2_2
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05589__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08070_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ net396 _03026_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ _03588_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05282_ _00994_ vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07021_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\] _00831_ net300 team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\]
+ _02675_ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05405__B2 _01069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08972_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] net827
+ net447 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__mux2_1
X_07923_ _03312_ _03477_ _03317_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__a21oi_1
Xhold18 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__A1 _02060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07028__C net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07854_ _03364_ _03389_ _03402_ _03403_ _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__o221a_1
X_06805_ _02466_ _02467_ _02468_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__or3_1
X_07785_ _01115_ net112 vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__nor2_1
X_04997_ net35 net34 net37 net36 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__or4_1
X_09524_ _00665_ _00666_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__nor2_1
X_06736_ _02406_ _02407_ _02408_ _02326_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recHEART.heartDetect
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_78_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10459__Q team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[3\]
+ net272 _04599_ net290 net220 vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a221o_1
X_06667_ _02108_ _02312_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__nor2_1
X_08406_ _03709_ _03880_ _03742_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__o21a_1
X_05618_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] _01327_
+ _01330_ _01324_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09386_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ _01424_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__nor2_1
X_06598_ net254 _02270_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__nor2_2
X_08337_ _03715_ _03813_ _03752_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_117_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05549_ _01259_ _01261_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08268_ _03709_ _03746_ _03742_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07219_ _02856_ _02860_ _01744_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08199_ net461 _01255_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__nand2_1
X_10230_ clknet_leaf_82_wb_clk_i _00041_ net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ clknet_leaf_3_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[8\]
+ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10092_ clknet_leaf_31_wb_clk_i team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[1\]
+ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_22_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05962__B _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10994_ net635 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_97_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10861__537 vssd1 vssd1 vccd1 vccd1 _10861__537/HI net537 sky130_fd_sc_hd__conb_1
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07085__B1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10428_ clknet_leaf_13_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[2\]
+ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06045__D1 _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10359_ clknet_leaf_23_wb_clk_i net726 net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.rand_num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06033__B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06060__A1 _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04920_ net3 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_109_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06036__D_N _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ _02208_ _03126_ _03127_ _03128_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06521_ _02088_ _02194_ _01646_ _01739_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09240_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ _04444_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06452_ _02125_ _02123_ _02122_ _02121_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__and4b_1
XFILLER_0_8_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05403_ net194 _01025_ _01102_ _01068_ _01038_ vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__o32a_1
X_09171_ net210 _04393_ _04394_ net402 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__a32o_1
XFILLER_0_111_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06383_ _01675_ _02056_ _02054_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__o21a_1
X_08122_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ _03608_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__or2_1
X_05334_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ _01046_ vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__and2_1
XANTENNA__06418__A3 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ net451 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ net393 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05265_ _00975_ _00977_ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout112_A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07004_ _00713_ _02666_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__xnor2_1
X_05196_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00904_ vssd1 vssd1
+ vccd1 vccd1 _00909_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06224__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ net476 _00827_ _01431_ _04244_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_129_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout481_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07906_ _03373_ _03459_ _03460_ _03457_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a31o_1
X_08886_ net439 _04208_ vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08879__A1 _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07837_ _03288_ _03351_ _03390_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__nand3b_1
XANTENNA__07551__A1 _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07551__B2 _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ _01083_ net186 vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__nor2_1
X_09507_ net869 net206 _04631_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06719_ _02390_ _02391_ _02389_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07699_ net108 _03253_ _03254_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__or3_1
XFILLER_0_91_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09438_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ _01415_ _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09369_ net226 _04535_ _04536_ net409 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05022__B _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05617__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05957__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10213_ clknet_leaf_81_wb_clk_i _00217_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_37_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input42_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05973__A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ clknet_leaf_1_wb_clk_i net721 net308 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_118_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10075_ clknet_leaf_35_wb_clk_i _00133_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07542__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06345__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06750__C1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10977_ net618 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_100_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05867__B net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold307 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[16\]
+ vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\] vssd1 vssd1
+ vccd1 vccd1 net988 sky130_fd_sc_hd__dlygate4sd3_1
X_05050_ _00776_ _00775_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold329 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05883__A _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08740_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ net239 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__mux2_1
X_05952_ net181 _01645_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__nor2_4
XANTENNA__06050__Y _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08671_ _04096_ _04097_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__a21o_1
X_05883_ _01574_ _01575_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_124_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07622_ _03119_ _03179_ _03176_ _03170_ _03168_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_124_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07553_ _01660_ _03080_ _03111_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__a21oi_1
X_10948__589 vssd1 vssd1 vccd1 vccd1 _10948__589/HI net589 sky130_fd_sc_hd__conb_1
XFILLER_0_76_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06504_ _02148_ _02176_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__nand2_4
X_07484_ _02278_ _03042_ _03043_ _01659_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09223_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ _04430_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__or2_1
XANTENNA__05123__A team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06435_ net279 _00753_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__and2_4
XFILLER_0_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout327_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07049__B1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04379_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__or2_1
X_06366_ net106 _01698_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__nor2_4
X_08105_ net753 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_cs _00244_
+ vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__o21ai_1
X_05317_ net191 _01004_ _01014_ vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ _04328_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06297_ net438 _01396_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout115_X net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06225__Y _01905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06272__A1 _00684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08036_ _03570_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ net393 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05248_ net492 _00797_ _00960_ vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__or3_2
XFILLER_0_101_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05179_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00886_ vssd1 vssd1
+ vccd1 vccd1 _00892_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09987_ clknet_leaf_45_wb_clk_i net415 net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07772__B2 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\] _04234_
+ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__and2_1
XANTENNA__07509__D1 _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06401__B _02060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ net264 _04192_ _04197_ _04195_ vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900_ net566 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_4_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07072__X _02726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10831_ net507 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_15_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07232__B _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10762_ clknet_leaf_66_wb_clk_i _00583_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10693_ clknet_leaf_70_wb_clk_i _00524_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05968__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06263__A1 _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10359__RESET_B net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07212__B1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08960__A0 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ clknet_leaf_36_wb_clk_i _00165_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_10058_ clknet_leaf_35_wb_clk_i net748 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07515__A1 _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910__655 vssd1 vssd1 vccd1 vccd1 net655 _10910__655/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_102_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10867__543 vssd1 vssd1 vccd1 vccd1 _10867__543/HI net543 sky130_fd_sc_hd__conb_1
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_69_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06039__A net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06220_ _01868_ _01871_ _01854_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06151_ net96 _01831_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__nand2_1
XANTENNA__07046__A3 _02699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05102_ net482 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\]
+ _00822_ _00824_ net1015 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__a32o_1
Xhold104 _00114_ vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold115 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[10\]
+ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06082_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] _01766_ _01761_
+ _01748_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__o211a_1
Xhold126 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09910_ _01780_ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__nand2_1
X_05033_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[0\]
+ _00764_ vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__o21ai_1
Xhold159 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09841_ _00657_ _04848_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06061__X _01748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06502__A _01582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[4\] vssd1 vssd1 vccd1 vccd1
+ _04797_ sky130_fd_sc_hd__nand3_1
X_06984_ _00712_ _00714_ _02645_ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__or3b_1
XANTENNA__06221__B net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08723_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[0\]
+ _04034_ _04082_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__a31o_1
X_05935_ net119 net111 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout277_A _00752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08654_ _04079_ _04081_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05866_ _01552_ _01556_ _01553_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__a21oi_1
X_07605_ net156 net107 _03161_ _03163_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__a31o_1
X_08585_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[20\]
+ _03622_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05797_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\] _01485_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] vssd1 vssd1
+ vccd1 vccd1 _01491_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07536_ _02223_ _03093_ _03094_ _01612_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_49_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07467_ net413 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ net395 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10439__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06418_ net107 net141 net166 _02091_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__a31o_2
XANTENNA__06493__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07690__B1 _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07398_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\] _02990_
+ net484 vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09137_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06349_ net418 net134 _02016_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__o31a_1
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05300__B _01005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09068_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08019_ net56 net40 net42 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__and3b_1
XFILLER_0_103_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout92_A _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08103__S _02671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06131__B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06181__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08058__B net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06720__A2 _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10814_ clknet_leaf_32_wb_clk_i team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.playButtonPixel
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08458__C1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08773__S net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10745_ clknet_leaf_67_wb_clk_i _00575_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10676_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[8\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06236__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06787__A2 _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07984__A1 _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07200__A3 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06041__B _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05720_ net1041 _00824_ _00825_ net1065 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05651_ _01352_ _01354_ _01357_ _01363_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06711__A2 _02262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08370_ net488 _00727_ _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__and3_1
X_05582_ _01286_ _01292_ _01294_ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__and3b_1
XFILLER_0_85_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07321_ net429 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07252_ _02898_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[5\]
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_119_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06203_ net94 _01879_ _01880_ net110 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07183_ net163 _01699_ _01718_ _01829_ net205 vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__o311a_1
XFILLER_0_121_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06134_ _01812_ _01813_ net285 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06065_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05016_ net288 net287 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__nand2_1
Xfanout403 net405 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_2
Xfanout414 net415 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout425 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\] vssd1
+ vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07727__A1 _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[2\] vssd1 vssd1
+ vccd1 vccd1 net436 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09824_ _04827_ _04836_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__nor2_1
XANTENNA__07047__B net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout447 net448 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_4
Xfanout458 team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1 vssd1 vccd1
+ vccd1 net458 sky130_fd_sc_hd__buf_2
Xfanout469 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[3\] vssd1
+ vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_2
X_09755_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\] _04783_ vssd1
+ vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__and2_1
X_06967_ net105 _02497_ _02543_ _02627_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout182_X net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06950__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05918_ net100 net87 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__or2_1
X_08706_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ _04121_ _04124_ _04115_ vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__o22a_1
X_09686_ net1107 _04735_ _04737_ _04730_ _04734_ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__o221a_1
X_06898_ net274 _02568_ _02562_ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_96_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08637_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ _04064_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__xnor2_1
X_10963__604 vssd1 vssd1 vccd1 vccd1 _10963__604/HI net604 sky130_fd_sc_hd__conb_1
X_05849_ _01538_ _01542_ _01536_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_7_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08568_ net54 net52 net139 vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__and3b_1
XFILLER_0_7_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07519_ _01873_ _02744_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__nor2_1
X_08499_ _03964_ _03965_ vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10530_ clknet_leaf_25_wb_clk_i _00398_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout87 _01610_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_4
XFILLER_0_107_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout98 net99 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06407__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10461_ clknet_leaf_22_wb_clk_i net1022 net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_91_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10392_ clknet_leaf_11_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[2\]
+ net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout95_X net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07238__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11013_ net390 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08768__S net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10754__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10728_ clknet_leaf_79_wb_clk_i _00558_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ clknet_leaf_3_wb_clk_i _00514_ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload13 clknet_leaf_89_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__inv_12
XFILLER_0_113_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload24 clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__inv_6
Xclkload35 clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_51_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload46 clknet_leaf_72_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__inv_6
XANTENNA__06209__B2 _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload57 clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_114_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload68 clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_114_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload79 clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__05875__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06052__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__B1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916__661 vssd1 vssd1 vccd1 vccd1 net661 _10916__661/LO sky130_fd_sc_hd__conb_1
X_07870_ _03361_ _03424_ _03419_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07185__A2 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ net90 _02467_ _02474_ _02491_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__o31ai_1
Xclkbuf_leaf_84_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09540_ _01419_ net291 _04645_ net270 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[37\]
+ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__a32o_1
X_06752_ net429 _00981_ net182 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09331__B1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05703_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ _01415_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_13_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07456__A_N net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09471_ net915 net207 _04608_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__o21a_1
X_06683_ _02345_ _02346_ _02355_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__and3_1
X_08422_ _03894_ _03896_ _03888_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__o21a_1
XANTENNA__05115__B net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05634_ net442 _01280_ _01327_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08353_ _03760_ _03825_ _03827_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__a31o_1
X_05565_ _01274_ _01277_ _01276_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__or3b_2
XANTENNA_fanout142_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07304_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08284_ net474 _03761_ _03760_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload7 clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_6
X_05496_ net422 _00690_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07235_ _02876_ _02879_ _02881_ _02885_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__o31a_1
XFILLER_0_73_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07660__A3 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07166_ _02799_ _02816_ _02818_ _02806_ _02814_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[1\]
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07948__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06117_ _01532_ _01797_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__nand2_2
XANTENNA__08070__B1 _03026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07097_ _02138_ net81 _02732_ _02750_ vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__a22o_1
XANTENNA__05959__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07058__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06048_ net163 _01735_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__nor2_2
Xfanout200 _01517_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_4
Xfanout211 _04376_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_2
Xfanout233 _02984_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_2
Xfanout244 net246 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_4
Xfanout255 net256 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07176__A2 _01901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 _00756_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_4
X_09807_ net247 vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__inv_2
Xfanout277 _00752_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05187__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout288 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[1\] vssd1
+ vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06384__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout299 _00969_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_4
X_07999_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__xor2_1
X_09738_ _04767_ _04771_ _04773_ net248 net1027 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__a32o_1
XFILLER_0_97_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09669_ _04716_ _04725_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_84_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07521__A _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06408__Y _02082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ clknet_leaf_18_wb_clk_i _00381_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05976__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10444_ clknet_leaf_39_wb_clk_i _00328_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07939__A1 _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10375_ clknet_leaf_12_wb_clk_i net694 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06611__A1 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06611__B2 _02282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06375__B1 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09313__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07150__B net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05350_ _01062_ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
XANTENNA__08961__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06047__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05281_ _00976_ _00978_ vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07020_ net398 _02674_ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06334__X _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06053__Y _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ net419 net792 net448 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__mux2_1
X_07922_ _01067_ net178 vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__nand2_1
Xhold19 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07853_ _03379_ _03404_ _03406_ _03407_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__or4_1
XANTENNA__06510__A _02135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ net90 _02474_ _02471_ net95 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_78_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07784_ _01058_ net108 vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nand2_1
X_04996_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[0\] vssd1 vssd1
+ vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06735_ _02311_ _02356_ _01413_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09523_ net922 net206 _04639_ vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout357_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09454_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ _04598_ _04597_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06666_ net99 _01616_ _02312_ net278 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_8_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08405_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03879_ _00727_
+ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__o21a_1
X_05617_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] _01319_
+ _01325_ _01315_ _01329_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__o221a_1
X_09385_ _00659_ _04546_ _04547_ _04542_ vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06597_ net158 _02021_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout145_X net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ net465 _03803_ _03812_ _03797_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o22a_1
X_05548_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] vssd1 vssd1 vccd1
+ vccd1 _01261_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08871__S net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08291__B1 _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ net416 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03745_
+ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05479_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_cleared _01191_ vssd1 vssd1
+ vccd1 vccd1 _01192_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07633__A3 _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07218_ _01645_ _01734_ _02867_ _02868_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06244__X _01921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08198_ net461 _01379_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07149_ _02800_ _02801_ _02798_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__o21a_1
X_10160_ clknet_leaf_3_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[7\]
+ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10091_ clknet_leaf_31_wb_clk_i team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[0\]
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09543__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10969__610 vssd1 vssd1 vccd1 vccd1 _10969__610/HI net610 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10993_ net634 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_57_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07085__A1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902__568 vssd1 vssd1 vccd1 vccd1 _10902__568/HI net568 sky130_fd_sc_hd__conb_1
XFILLER_0_34_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10427_ clknet_leaf_13_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[1\]
+ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06045__C1 _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ clknet_leaf_6_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear
+ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.maze_clear_edge_detector.inter
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10289_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[2\]
+ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_109_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06899__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06520_ net205 _02089_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__or2_2
XFILLER_0_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06451_ net168 _01711_ _01734_ _02058_ _02092_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06048__Y _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05402_ net397 _01058_ vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__nand2_2
X_09170_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04391_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06382_ net181 _01873_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__or2_4
X_08121_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[3\]
+ _03607_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05333_ _00966_ net299 _01045_ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08052_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ net298 _03579_ vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05264_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ _00973_ vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07003_ _02649_ _02665_ _02648_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_40_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05195_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00901_ vssd1 vssd1
+ vccd1 vccd1 _00908_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout105_A _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08954_ net492 _00797_ _01427_ _01428_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_129_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07905_ net259 _03382_ _03385_ _03386_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__nor4_1
X_08885_ _04205_ _04207_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__or2_1
X_07836_ _03390_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__inv_2
XANTENNA__07551__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04979_ net474 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ _01084_ net189 vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09506_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[23\]
+ net271 net292 net222 vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__a211o_1
X_06718_ _02066_ _02313_ net83 net253 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a22oi_1
X_07698_ net278 net93 net115 net88 _02009_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06649_ _02127_ _02297_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__nand2_1
X_09437_ net417 _01414_ _04585_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09368_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04533_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07067__B2 _02110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ net415 net465 vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09299_ net963 net404 net229 _04487_ vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06814__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10212_ clknet_leaf_83_wb_clk_i _00216_ net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_37_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10143_ clknet_leaf_1_wb_clk_i net734 net308 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05973__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819__495 vssd1 vssd1 vccd1 vccd1 _10819__495/HI net495 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_89_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input35_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ clknet_leaf_34_wb_clk_i _00132_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07542__A2 _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08077__A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10976_ net617 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_58_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05988__X _01681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06325__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold308 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\] vssd1 vssd1 vccd1
+ vccd1 net978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold319 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[19\]
+ vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06281__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06569__B1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07230__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05883__B _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05951_ net184 net176 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__nand2_8
X_08670_ _04054_ _04058_ _04073_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__a31o_1
X_05882_ _01574_ _01575_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_124_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07621_ _03177_ _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_124_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07552_ _01739_ net165 _03110_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06503_ _02148_ _02176_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_17_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07483_ _02278_ _03042_ _03043_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09222_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ _04430_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__nand2_1
X_06434_ net267 _02030_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__or2_4
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08715__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09153_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ _04379_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__nand2_1
XANTENNA__07049__A1 _01921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06365_ _02034_ _02035_ _02038_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__and3_1
XANTENNA__07049__B2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08104_ net789 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataDc _02671_
+ vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__mux2_1
X_05316_ _01026_ _01028_ vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__or2_1
X_09084_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ _04328_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__nand2_1
X_06296_ net162 _01969_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08035_ net413 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net294 _03569_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a221o_1
X_05247_ _00683_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_cleared vssd1
+ vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__or2_4
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout108_X net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05178_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00890_ vssd1 vssd1
+ vccd1 vccd1 _00891_ sky130_fd_sc_hd__xnor2_1
X_09986_ clknet_leaf_86_wb_clk_i _00091_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07066__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ _01432_ _01484_ _01762_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__C1 _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10658__RESET_B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08868_ _00942_ _04196_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07819_ _01057_ net173 vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_84_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08799_ _04153_ _04154_ net196 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10830_ net506 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_95_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05314__A _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ clknet_leaf_67_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[8\]
+ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10692_ clknet_leaf_70_wb_clk_i _00523_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05968__B net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05984__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06432__X _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07212__A1 _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ clknet_leaf_27_wb_clk_i _00164_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05990__Y _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ clknet_leaf_29_wb_clk_i net766 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07515__A2 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07704__A _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload0_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05224__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10959_ net600 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XFILLER_0_58_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10908__574 vssd1 vssd1 vccd1 vccd1 _10908__574/HI net574 sky130_fd_sc_hd__conb_1
XFILLER_0_6_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_38_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05230__Y _00943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06150_ net185 net176 _01657_ net102 _01830_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__a41o_1
XFILLER_0_108_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06055__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05101_ net481 team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00810_ _00816_
+ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__and4_2
XFILLER_0_124_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06081_ _01762_ _01767_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold105 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[7\] vssd1
+ vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold138 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_num\[0\]
+ vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__dlygate4sd3_1
X_05032_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__nor2_1
Xhold149 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08270__A _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09840_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\] _04844_ vssd1
+ vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__and2_1
XANTENNA__05214__B1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06502__B net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09771_ _04796_ _04794_ net997 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__mux2_1
X_06983_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\] _02645_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] vssd1 vssd1
+ vccd1 vccd1 _02647_ sky130_fd_sc_hd__a21o_1
X_08722_ _04135_ _04134_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__mux2_1
X_05934_ net117 _01616_ _01626_ net87 net101 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__a311oi_4
XANTENNA__09900__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08653_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01239_ _04080_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__or3_1
X_05865_ _01547_ net158 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07604_ net137 _01688_ _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__and3_1
X_08584_ net146 _04026_ _03965_ vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__a21o_1
XANTENNA__06190__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05796_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] _01486_
+ _01487_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07535_ net100 _02107_ _02191_ _03072_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout437_A team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07466_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ net294 _03034_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[28\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06517__X _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09205_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06417_ net216 net175 _01698_ _01684_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06493__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07397_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\] _02990_
+ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__and2_1
XANTENNA__07690__B2 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06348_ _02012_ _02022_ _02019_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__or3b_1
X_09136_ net4 net1181 _04368_ vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09067_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ net6 _04317_ vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06279_ net204 _01954_ _01955_ _01952_ _01944_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08018_ net1070 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_back
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05205__B1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ clknet_leaf_83_wb_clk_i _00074_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_51_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06131__C _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07524__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10813_ clknet_leaf_78_wb_clk_i _00634_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08458__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10744_ clknet_leaf_72_wb_clk_i _00574_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07130__B1 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10675_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[7\]
+ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08642__X _04070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05985__Y _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07984__A2 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10834__510 vssd1 vssd1 vccd1 vccd1 _10834__510/HI net510 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_8_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10109_ clknet_leaf_55_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireHighlightDetect
+ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05650_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] _01301_
+ _01362_ _01360_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08964__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05581_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] _01253_
+ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07320_ _01190_ _01192_ _01193_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07251_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ _02897_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07672__A1 _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07672__B2 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06202_ net110 _01880_ _01881_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07182_ _02134_ net82 _02741_ _02831_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06133_ _01812_ _01813_ net284 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08712__B net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07609__A _02254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06064_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06072__X _01759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05015_ _00649_ net280 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__nor2_4
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_2
XFILLER_0_100_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07188__B1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout415 _00017_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07727__A2 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout426 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_4
Xfanout437 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] vssd1 vssd1
+ vccd1 vccd1 net437 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09823_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\] _04834_ vssd1
+ vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__and2_1
Xfanout448 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.activate_rand_delay_2
+ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_4
Xfanout459 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\] vssd1 vssd1
+ vccd1 vccd1 net459 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout387_A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ net978 _04782_ _04784_ net248 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__o22a_1
X_06966_ _02488_ _02560_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__nand2_1
X_08705_ _04122_ _04123_ net243 vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07344__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05917_ net92 _01609_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__nand2_1
X_09685_ _04730_ _04737_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout175_X net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06897_ _02549_ _02567_ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ _00693_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__or2_1
XANTENNA__06163__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05848_ _01540_ _01541_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08567_ _03615_ _04014_ net139 vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a21oi_1
X_05779_ _01468_ _01471_ _01473_ _01459_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_7_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07518_ net184 _01657_ net260 vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__a21oi_2
X_08498_ _02670_ _03626_ _03652_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__nor3_2
XFILLER_0_9_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07449_ net453 net451 vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__and2_2
Xfanout88 _01609_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout99 _01600_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06407__B _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10460_ clknet_leaf_13_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_down
+ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09119_ net212 _04354_ _04356_ net399 net1035 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__a32o_1
X_10391_ clknet_leaf_11_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[1\]
+ net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06423__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10673__RESET_B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07238__B _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold480 team_07_WB.instance_to_wrap.team_07.label_num_bus\[24\] vssd1 vssd1 vccd1
+ vccd1 net1150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold491 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout88_X net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ net640 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_99_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05981__B _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07639__D1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10727_ clknet_leaf_79_wb_clk_i _00557_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07654__A1 _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05221__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10658_ clknet_leaf_3_wb_clk_i _00513_ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkload14 clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__inv_6
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload25 clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_113_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload36 clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__08603__B1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload47 clknet_leaf_74_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10589_ clknet_leaf_37_wb_clk_i _00453_ net363 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload58 clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__inv_8
XFILLER_0_11_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06604__Y _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload69 clknet_leaf_38_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_114_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08959__S _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06052__B net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__A2 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ net89 _02467_ _02477_ net111 _02490_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__a221o_1
X_10986__627 vssd1 vssd1 vccd1 vccd1 _10986__627/HI net627 sky130_fd_sc_hd__conb_1
X_06751_ net429 _00981_ net182 _02420_ _02422_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a32o_1
X_05702_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\] vssd1
+ vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__or2_2
X_06682_ _02336_ _02339_ _02343_ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__or3b_1
X_09470_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[10\]
+ net273 net292 net222 vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__a211o_1
XANTENNA__06145__B2 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07451__X _03026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08421_ _03656_ _03667_ _03895_ _03890_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05633_ net442 _01322_ _01344_ _01345_ _01320_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08352_ _03760_ _03825_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_53_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_05564_ _01266_ _01270_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07303_ net444 _01328_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08283_ net467 _03643_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__nand2_1
X_05495_ net422 _00690_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload8 clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__06227__B _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout135_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07234_ _02882_ _02884_ _02880_ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__or3b_1
XFILLER_0_41_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07165_ net168 _02033_ _02758_ _02817_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__a31o_1
XFILLER_0_125_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06116_ net177 net123 _01702_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__or3_2
X_07096_ _01618_ _01921_ _02196_ net265 _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__a221o_2
XANTENNA__06243__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05959__A1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06047_ net128 _01699_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__nand2_4
XFILLER_0_2_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07058__B _02209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10084__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout201 _01517_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_4
Xfanout212 _04325_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_2
Xfanout223 _04582_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_2
Xfanout234 net235 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_4
Xfanout245 net246 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_8
Xfanout256 net257 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_4
X_09806_ _04798_ _04804_ _04807_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__o21ai_2
Xfanout267 _00747_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_4
XANTENNA__09570__A1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__A2 _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 _00651_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_4
XANTENNA__06384__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout289 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[1\] vssd1
+ vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_2
X_07998_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__xor2_1
XANTENNA__07581__B1 _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ _04772_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__inv_2
X_06949_ net174 _02506_ _02508_ _02581_ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_69_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09668_ _04716_ _04724_ _04725_ vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__nor3_1
XANTENNA__07333__A0 _00675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08619_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ net457 vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__or2_1
X_09599_ _04665_ _04675_ net1113 vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07636__A1 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10512_ clknet_leaf_18_wb_clk_i _00380_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10443_ clknet_leaf_46_wb_clk_i net811 net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07939__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10374_ clknet_leaf_11_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[2\]
+ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06611__A2 _02073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05992__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__X _03095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06375__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05216__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09864__A2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08824__B1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06047__B _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05280_ _00988_ _00992_ vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__nand2_2
XFILLER_0_102_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10595__RESET_B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05886__B _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08970_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] net785
+ net448 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__mux2_1
X_07921_ net131 net122 _03475_ _03473_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__a31o_1
X_07852_ net105 _03376_ _03387_ net106 vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06510__B _02178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06803_ net434 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1 vssd1
+ vccd1 vccd1 _02474_ sky130_fd_sc_hd__xnor2_2
Xinput1 gpio_in[22] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_1
X_07783_ _03285_ _03286_ _03337_ _03336_ _03335_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__o32a_1
XANTENNA__06563__A1_N _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04995_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\] vssd1 vssd1
+ vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
XANTENNA__08107__A2 _02671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[31\]
+ net270 _04638_ net223 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a211o_1
X_06734_ _02307_ _02359_ _01223_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09453_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\] vssd1
+ vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__and2b_1
X_06665_ _02334_ _02336_ _02337_ _02330_ _02259_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__o32a_1
XFILLER_0_66_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08404_ _03745_ _03804_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__nor2_1
X_05616_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] net444
+ _01328_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__a21o_1
X_09384_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[16\]
+ net409 _04308_ net226 vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__a22o_1
X_06596_ _02267_ _02264_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08335_ _03718_ _03811_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__nor2_1
X_05547_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout138_X net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07094__A2 _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05478_ _00795_ _00963_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__o21ai_1
X_08266_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\] _03744_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07633__A4 _03117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07217_ net183 _02033_ _02863_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08197_ net460 _01381_ _03675_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07148_ _02072_ _02758_ _02781_ _02059_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07079_ _02732_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__inv_2
X_10090_ clknet_leaf_68_wb_clk_i _00148_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06701__A _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10992_ net633 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06148__A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05987__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07085__A2 _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06435__X _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10426_ clknet_leaf_13_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[0\]
+ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06045__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10357_ clknet_leaf_59_wb_clk_i _00297_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10288_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[1\]
+ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07848__A1 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07848__B2 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06450_ net169 _01734_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__nand2_1
XANTENNA__08972__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06058__A _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10776__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05401_ _00970_ _01031_ _01089_ _01090_ _01101_ vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__o221a_1
X_06381_ net181 _01873_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__nor2_2
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08120_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[2\]
+ _03606_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__or2_1
X_05332_ _01018_ _01039_ _01044_ _01032_ vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__or4b_1
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08273__A _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08051_ net452 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ net394 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__a22o_1
X_05263_ net429 net430 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07002_ _02649_ _02664_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__xnor2_1
X_05194_ _00902_ _00903_ _00905_ _00906_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08953_ net490 _04243_ vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08328__A2 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07904_ net158 _03374_ _03458_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__or3b_1
X_08884_ _01399_ _01397_ _04203_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07835_ net278 _01055_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__nand2_1
X_07766_ _03307_ _03319_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__nor2_1
X_04978_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.cs vssd1 vssd1 vccd1
+ vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_cs sky130_fd_sc_hd__inv_2
XFILLER_0_56_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09505_ net886 net222 _04605_ net920 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06717_ _02079_ _02258_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07697_ net119 _02031_ _02148_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__o21ai_1
X_09436_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\] vssd1
+ vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__and2b_1
X_06648_ _02080_ _02287_ _02289_ _02135_ _02320_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04533_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__or2_1
X_06579_ _01627_ _02106_ _02149_ _02251_ _02252_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10999__637 vssd1 vssd1 vccd1 vccd1 _10999__637/HI net637 sky130_fd_sc_hd__conb_1
XANTENNA__10446__RESET_B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08318_ _03722_ _03795_ _03718_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_10_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09298_ _04485_ _04486_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05078__B2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06814__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ net462 _01282_ _01308_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06415__B _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10211_ clknet_leaf_81_wb_clk_i _00215_ net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_37_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10142_ clknet_leaf_1_wb_clk_i _00042_ net308 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_37_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10073_ clknet_leaf_35_wb_clk_i _00131_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07527__B1 _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06750__A1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10975_ net616 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_43_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06606__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold309 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[10\]
+ vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ clknet_leaf_14_wb_clk_i _00300_ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[2\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07230__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06341__A _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05950_ net188 net173 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__nor2_1
XANTENNA__08967__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07518__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05881_ _01565_ _01573_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__or2_4
XANTENNA__08191__B1 _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07620_ _01721_ _03079_ _03120_ _01733_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_124_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07613__A2_N net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07551_ _01658_ net172 _01701_ _01669_ _01664_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__o32a_1
XFILLER_0_88_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06502_ _01582_ net115 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_17_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07482_ net255 net187 _01901_ _01664_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09221_ net230 _04431_ _04432_ net406 net890 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__a32o_1
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06433_ net267 _02030_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__nor2_4
XFILLER_0_91_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08274__Y _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09152_ net210 _04380_ _04381_ net399 net941 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06364_ _01685_ _02036_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08103_ net778 _03604_ _02671_ vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05315_ net194 _01027_ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__nor2_1
X_06295_ net148 _01966_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__or2_1
X_09083_ net213 _04329_ _04330_ net400 net912 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout215_A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ net454 net451 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__and3_1
X_05246_ _00957_ _00958_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05177_ _00888_ _00889_ _00873_ vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__mux2_2
X_09985_ clknet_leaf_81_wb_clk_i _00090_ net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851__527 vssd1 vssd1 vccd1 vccd1 _10851__527/HI net527 sky130_fd_sc_hd__conb_1
XANTENNA__07066__B _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] net1141 net241 vssd1
+ vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08867_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] _00941_ vssd1 vssd1
+ vccd1 vccd1 _04196_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07818_ _01058_ net179 vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_84_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08798_ net341 _01450_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07749_ _01084_ _01566_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10760_ clknet_leaf_67_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[7\]
+ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09419_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\] _04567_
+ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__nand3_1
XANTENNA__07810__A _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05463__A2_N _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10691_ clknet_leaf_53_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[23\]
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06799__A1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05984__B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07212__A2 _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10312__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ clknet_leaf_27_wb_clk_i _00163_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10056_ clknet_leaf_35_wb_clk_i net774 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10368__RESET_B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05224__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10958_ net599 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_70_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06487__B1 _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07720__A _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10889_ net646 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_26_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08027__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08779__A2 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10407__SET_B net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06055__B net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05100_ net1041 _00817_ _00823_ net1016 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06080_ _00655_ _01766_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold106 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07014__A_N team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.idle vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold117 _00110_ vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__dlygate4sd3_1
X_05031_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _00762_ vssd1
+ vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold139 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_78_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10954__595 vssd1 vssd1 vccd1 vccd1 _10954__595/HI net595 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\] _04767_ _04790_
+ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__and3_1
X_06982_ _00714_ _02645_ vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08721_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _04134_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__nor2_1
X_05933_ net276 _01625_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08652_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.wait_cnt\[0\]
+ _04071_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_1_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05864_ _01548_ _01550_ _01551_ _01555_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_1_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06714__A1 _02135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ _03063_ _03093_ _03072_ _02182_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a2bb2o_1
X_08583_ _03621_ _04025_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__nand2_1
X_05795_ _01486_ _01487_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__nand2_1
XANTENNA__06190__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07534_ _02779_ _03092_ _01619_ _02119_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06478__B1 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07465_ net413 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ net396 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout332_A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06416_ _02087_ _02088_ _02089_ _01711_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06493__A3 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07396_ _02990_ _02991_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[4\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07690__A2 _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06246__A team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09135_ _04321_ _04364_ _04365_ _04367_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__or4_1
X_06347_ _02018_ _02020_ _02021_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout120_X net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout218_X net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09066_ _04307_ _04309_ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06278_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] _01941_ _01948_ vssd1
+ vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_115_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05453__A1 _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ net1044 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_select
+ sky130_fd_sc_hd__and2b_1
X_05229_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] _00941_ vssd1 vssd1
+ vccd1 vccd1 _00942_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10892__649 vssd1 vssd1 vccd1 vccd1 net649 _10892__649/LO sky130_fd_sc_hd__conb_1
XANTENNA__07077__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ clknet_leaf_87_wb_clk_i _00073_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_51_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08919_ _04222_ _04223_ _04225_ _04227_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__or4b_2
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09899_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\] _01777_
+ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07524__B _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06705__A1 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06181__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10812_ clknet_leaf_78_wb_clk_i _00633_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07540__A _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10743_ clknet_leaf_72_wb_clk_i _00573_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07130__A1 _01694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10674_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[6\]
+ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07969__B1 _01681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07539__X _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05995__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07197__A1 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07197__B2 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05219__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10108_ clknet_leaf_55_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[5\]
+ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10039_ _00059_ _00637_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06172__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05580_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] _01253_
+ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07250_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07672__A2 _02055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06201_ _01881_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07181_ _02138_ net81 _02750_ _02831_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07449__X _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06132_ net127 _01699_ net158 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06063_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05014_ net268 net267 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__nand2_1
XANTENNA__07188__A1 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout405 net410 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_2
Xfanout416 team_07_WB.instance_to_wrap.team_07.heartPixel vssd1 vssd1 vccd1 vccd1
+ net416 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09822_ _04827_ _04834_ _04835_ vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__nor3_1
Xfanout427 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_4
XFILLER_0_39_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout438 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[2\] vssd1 vssd1 vccd1
+ vccd1 net438 sky130_fd_sc_hd__buf_2
Xfanout449 net450 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_4
X_09753_ _00652_ _04783_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__nor2_1
X_06965_ _02602_ _02634_ _02635_ net268 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout282_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _01238_ _04062_ _01240_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__a21o_1
X_05916_ _01582_ _01597_ _01604_ net120 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__and4_2
X_09684_ _04736_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__inv_2
X_06896_ _02564_ _02565_ _02566_ _02486_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__or4b_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10219__RESET_B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06699__B1 _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08635_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ _04062_ net457 vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__o21ai_1
X_05847_ _01508_ _01519_ _01539_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout168_X net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08566_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[12\]
+ _03614_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05371__B1 _01067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05778_ net414 _01476_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__nor2_1
XANTENNA__05910__A2 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07517_ _03075_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08497_ net53 net146 _03959_ net1089 vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07112__A1 _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout335_X net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07448_ team_07_WB.EN_VAL_REG net392 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__or2_1
XFILLER_0_9_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout89 _01606_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05674__A1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06871__B1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07379_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\] _02979_
+ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09118_ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__inv_2
X_10390_ clknet_leaf_10_wb_clk_i net689 net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07966__A3 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09049_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ _04301_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__or2_1
X_10857__533 vssd1 vssd1 vccd1 vccd1 _10857__533/HI net533 sky130_fd_sc_hd__conb_1
XANTENNA__07519__B _02744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06423__B _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold470 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold481 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] vssd1 vssd1 vccd1
+ vccd1 net1151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 team_07_WB.instance_to_wrap.team_07.label_num_bus\[8\] vssd1 vssd1 vccd1
+ vccd1 net1162 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net390 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ clknet_leaf_79_wb_clk_i _00556_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05996__Y _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10657_ clknet_leaf_2_wb_clk_i _00512_ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload15 clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__clkinv_8
Xclkload26 clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_6
Xclkload37 clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10588_ clknet_leaf_37_wb_clk_i _00452_ net363 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.ssdec_sck
+ sky130_fd_sc_hd__dfrtp_1
Xclkload48 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__inv_8
XFILLER_0_50_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload59 clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_114_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06668__A2_N _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07709__A3 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_58 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06750_ net174 _02418_ _02421_ _00971_ net138 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__a221o_1
XANTENNA__08975__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05701_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\] vssd1
+ vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__nor2_1
XANTENNA__09331__A2 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06681_ _02351_ _02353_ _02327_ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08420_ net475 _03642_ _03665_ net469 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__o211ai_1
X_05632_ net442 _01327_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__nor2_1
XANTENNA__06696__A3 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05252__X _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08351_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\] _03826_
+ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05563_ _01273_ _01275_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07302_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ _02925_ _02928_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[5\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08282_ _00717_ _03643_ net467 vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__a21o_1
X_05494_ _01204_ _01206_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload9 clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_8
XANTENNA__06227__C _01905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07233_ net129 _02773_ _02883_ _02874_ _02767_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__a32o_1
XFILLER_0_15_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_22_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07164_ net107 _01710_ _02761_ _02781_ _02803_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__a32o_1
XANTENNA__06524__A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06115_ net126 _01701_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08070__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07095_ _02109_ _02139_ _02735_ vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__o21a_1
XANTENNA__06243__B net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05959__A2 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06046_ net123 _01700_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__nor2_2
XFILLER_0_100_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout202 net203 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_4
Xfanout213 _04325_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_2
Xfanout224 net225 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_4
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_2
Xfanout246 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.activate_rand
+ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input2_A gpio_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _04823_ _04821_ net1042 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__mux2_1
Xfanout257 _01489_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_6
Xfanout268 _00746_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_4
X_07997_ _03548_ _03549_ vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__xnor2_1
Xfanout279 _00651_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07581__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06384__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__and4_1
X_06948_ _02615_ _02616_ _02618_ _02614_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__or4b_1
XFILLER_0_69_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09667_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[6\]
+ _04721_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06879_ _02543_ _02529_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__and2b_1
XFILLER_0_96_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08618_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ net457 vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__nor2_1
X_09598_ _04666_ _04674_ _04676_ _04664_ net1040 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__a32o_1
XFILLER_0_55_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07090__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10928__578 vssd1 vssd1 vccd1 vccd1 _10928__578/HI net578 sky130_fd_sc_hd__conb_1
X_08549_ net1160 _03610_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10511_ clknet_leaf_18_wb_clk_i _00379_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ clknet_leaf_46_wb_clk_i _00326_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_94_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06434__A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10373_ clknet_leaf_11_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[1\]
+ net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05992__B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06375__A2 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06609__A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07875__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ clknet_leaf_71_wb_clk_i _00540_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08052__A2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07920_ _03306_ _03445_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05247__X _00960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ net161 _03366_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__nor2_1
XANTENNA__08760__A0 team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06802_ net99 _02470_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__nand2_1
Xinput2 gpio_in[23] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_2
X_07782_ _01105_ _02212_ _02191_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__a21oi_1
X_04994_ net461 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09521_ _00665_ _01419_ net291 _04637_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__o211a_1
X_06733_ net424 net423 _02360_ _02361_ _02405_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__a311o_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09452_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\] net417
+ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__o21ai_1
X_06664_ _01626_ _02258_ _01638_ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08403_ _03858_ _03877_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__or2_1
X_05615_ net445 net443 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__or2_1
X_09383_ net226 _04545_ _04546_ net408 net932 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__a32o_1
X_06595_ net262 _02264_ _02265_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout245_A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05142__B team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08334_ _03809_ _03810_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05546_ net421 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] vssd1 vssd1 vccd1
+ vccd1 _01259_ sky130_fd_sc_hd__or3_2
XFILLER_0_74_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05629__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08265_ net4 _00660_ _00663_ _03704_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__a41o_2
XFILLER_0_117_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05477_ _01153_ _01174_ _01189_ _01046_ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08453__B _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07216_ _02065_ net82 _02736_ _02861_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08196_ _00678_ net460 _01254_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07147_ net104 _02277_ _02761_ net166 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout200_X net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07078_ _02726_ _02729_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06029_ net136 net128 net145 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__a21oi_4
XANTENNA_input5_X net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09719_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\]
+ _04754_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\] vssd1 vssd1
+ vccd1 vccd1 _04760_ sky130_fd_sc_hd__a31o_1
X_10991_ net632 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_87_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06148__B _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08644__A _04070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05987__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07490__B1 _03050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10425_ clknet_leaf_13_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[2\]
+ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10356_ clknet_leaf_57_wb_clk_i _00296_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10287_ clknet_leaf_44_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[0\]
+ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07545__B2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06339__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05400_ _01056_ _01094_ vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__nand2_2
XFILLER_0_28_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06380_ net202 net172 _01663_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__a21o_4
XFILLER_0_127_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05331_ _01035_ _01037_ _01043_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__or3b_1
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08050_ net1154 net298 _03578_ vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__a21o_1
X_05262_ _00673_ _00974_ vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07001_ _02664_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05193_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00904_ vssd1 vssd1
+ vccd1 vccd1 _00906_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06802__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08952_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_col
+ _04234_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared vssd1 vssd1
+ vccd1 vccd1 _04243_ sky130_fd_sc_hd__a31o_1
XANTENNA__05726__C_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08328__A3 _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ net134 _03366_ _03365_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__o21ba_1
X_08883_ _04206_ net1076 _04205_ vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout195_A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06240__C _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07834_ net106 _03380_ _03388_ _01692_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07765_ _03319_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_04977_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] vssd1
+ vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout362_A net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06716_ net144 _01737_ _02260_ _02388_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__a31o_1
X_09504_ net920 net206 _04630_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07696_ _01619_ net253 _02249_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__or3b_1
XFILLER_0_52_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09435_ _01429_ _01430_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__or2_2
X_06647_ _02067_ _02281_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout150_X net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09366_ net226 _04532_ _04534_ net409 net1123 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06578_ net283 net98 net119 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__and3_1
X_08317_ _03742_ _03794_ _03793_ net485 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__a211o_1
X_05529_ _01197_ _01240_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__nor2_1
X_09297_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ _04481_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08248_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] _03725_ _03726_
+ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08179_ _03644_ _03656_ _03657_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10415__RESET_B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10210_ clknet_leaf_83_wb_clk_i _00214_ net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ clknet_leaf_31_wb_clk_i team_07_WB.instance_to_wrap.team_07.recFLAG.flagDetect
+ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.flagPixel sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05786__B1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10072_ clknet_leaf_35_wb_clk_i _00130_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07527__A1 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05538__B1 _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07543__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10974_ net615 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XANTENNA__06159__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05998__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06606__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10408_ clknet_leaf_14_wb_clk_i _00299_ net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10339_ clknet_leaf_54_wb_clk_i _00279_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07230__A3 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07518__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05880_ _01569_ _01570_ _01572_ _01573_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__or4b_4
XFILLER_0_89_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07550_ net169 _02262_ _02219_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06501_ _02173_ _02174_ _02149_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07481_ _01658_ _01873_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09220_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a21o_1
X_06432_ net288 net286 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__or2_4
XFILLER_0_5_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09151_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06363_ net135 net126 net170 _01935_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__and4_1
XANTENNA__06075__Y _01762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ _03603_ _03602_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__mux2_1
XANTENNA__06516__B _02178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10959__600 vssd1 vssd1 vccd1 vccd1 _10959__600/HI net600 sky130_fd_sc_hd__conb_1
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05314_ _01010_ _01019_ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__or2_1
X_09082_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06294_ net148 _01966_ _01969_ net162 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_44_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08033_ _03568_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ net394 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__mux2_1
X_05245_ _00684_ _00946_ vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout208_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05176_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\]
+ _00883_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09984_ clknet_leaf_82_wb_clk_i _00089_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05148__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08935_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ net241 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__A1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07066__C net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout198_X net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ _00685_ _04192_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07817_ _01058_ net178 vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__nor2_1
X_08797_ net806 _04151_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07748_ _01068_ net159 vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07679_ _03161_ _03234_ _03236_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09418_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\]
+ _04572_ _04567_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__mux2_1
XANTENNA__07810__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10690_ clknet_leaf_53_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[22\]
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10667__RESET_B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09349_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ _04520_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06442__A _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10124_ clknet_leaf_29_wb_clk_i _00162_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input40_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10055_ clknet_leaf_35_wb_clk_i net763 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10957_ net598 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10888_ net645 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_26_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06336__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05571__C_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07987__B2 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold107 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold118 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[3\]
+ vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__dlygate4sd3_1
X_05030_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__or2_1
XANTENNA__07448__A team_07_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08043__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06352__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06981_ _02645_ _02646_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__nor2_1
X_08720_ _04034_ _04082_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__nand2_1
X_05932_ _01620_ _01625_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__and2_4
Xclkbuf_leaf_47_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08651_ _04066_ _04071_ _04078_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__and3_1
X_05863_ _01548_ _01550_ _01551_ _01555_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_1_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07602_ _03073_ _03160_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08582_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[18\]
+ _03620_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__nand2_1
X_05794_ _01486_ _01487_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07533_ _00759_ net99 net120 vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout158_A _01558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07464_ net453 net413 vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06527__A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09203_ net5 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ _04417_ vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__mux2_1
X_06415_ _01709_ _01720_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07395_ net1139 _02988_ net480 vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_33_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06246__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09134_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__or4_1
X_06346_ net177 _02014_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__or2_4
XFILLER_0_127_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07978__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09065_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04313_ _04315_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__nor4_1
XFILLER_0_130_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06277_ net458 net262 _01951_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout113_X net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08016_ net1021 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_right
+ sky130_fd_sc_hd__and2b_1
X_05228_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\] net450 vssd1 vssd1
+ vccd1 vccd1 _00941_ sky130_fd_sc_hd__nand2_1
XANTENNA__06650__A1 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05159_ _00865_ _00866_ _00871_ _00858_ vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__a31o_1
XANTENNA__07077__B net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ clknet_leaf_84_wb_clk_i _00072_ net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_08918_ _00724_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ _00725_ _04226_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__o221a_1
XANTENNA__07805__B net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ net855 net154 net151 _04886_ vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__a22o_1
XANTENNA__07093__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ net395 net393 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__o21a_1
XANTENNA__07524__C net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06705__A2 _02073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10413__SET_B net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811_ clknet_leaf_78_wb_clk_i _00632_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06469__B2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10742_ clknet_leaf_72_wb_clk_i _00572_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06437__A _02110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10673_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[5\]
+ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10430__RESET_B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07969__A1 _01113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05995__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07197__A2 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06900__A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10107_ clknet_leaf_55_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[4\]
+ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05462__D_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ _00058_ _00636_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10589__RESET_B net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06200_ _01863_ _01865_ _01864_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_30_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07180_ _02831_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10100__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06131_ net133 net121 _01677_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__or3_4
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06062_ _00687_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared _01238_
+ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__or3b_1
X_05013_ net267 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09582__A0 _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07188__A2 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout406 net407 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_2
X_09821_ _04825_ _04833_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__a21oi_1
Xfanout417 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[3\]
+ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_2
Xfanout428 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout439 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[2\] vssd1 vssd1 vccd1
+ vccd1 net439 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06810__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07184__Y _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[8\] _04777_ vssd1 vssd1
+ vccd1 vccd1 _04783_ sky130_fd_sc_hd__and4_1
X_06964_ _02487_ _02560_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08703_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _04067_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__or2_1
X_05915_ _01582_ net120 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__and2_2
X_09683_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[2\] vssd1 vssd1 vccd1
+ vccd1 _04736_ sky130_fd_sc_hd__and3_1
X_06895_ net115 _02476_ _02528_ _02539_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout275_A _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06699__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ _01196_ _04061_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__nand2_1
X_05846_ _01519_ _01539_ _01508_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07641__A _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08565_ _04012_ _04013_ _03996_ vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__o21a_1
X_05777_ _01475_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__inv_2
XANTENNA__05371__A1 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07516_ _02108_ _02150_ _03071_ _03073_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__o211a_1
X_08496_ net140 _03629_ _03960_ net54 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07112__A2 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07447_ net905 _03021_ _03023_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[23\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__06856__D1 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07378_ _02979_ _02980_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06329_ net123 _01963_ _01965_ _01993_ _01641_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a41o_1
X_09117_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ _04350_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09048_ _04301_ _04302_ net1121 net405 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold460 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07238__D _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout90_A _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold471 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net390 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
Xhold482 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[6\] vssd1
+ vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06387__B1 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06926__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05336__A team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06167__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10725_ clknet_leaf_79_wb_clk_i _00555_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10656_ clknet_leaf_2_wb_clk_i _00511_ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08382__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08064__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload16 clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_16
X_10587_ clknet_leaf_37_wb_clk_i _00451_ net363 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.ssdec_sdi
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload27 clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_134_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload38 clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__clkinv_8
Xclkload49 clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__inv_8
XFILLER_0_50_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09941__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05700_ net423 net425 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__nand2b_4
X_06680_ _00759_ _01627_ _02178_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__or3_1
XANTENNA__10325__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05631_ _01319_ _01343_ _00680_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__and3b_1
XANTENNA__10352__RESET_B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08350_ _03637_ _03815_ _03766_ _03632_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_47_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05562_ _01266_ _01274_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07301_ _02928_ _02929_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[4\]
+ sky130_fd_sc_hd__nor2_1
X_08281_ net469 _03756_ _03758_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05493_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ _01205_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06302__B1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07232_ _01936_ _02873_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__nor2_1
X_10923__668 vssd1 vssd1 vccd1 vccd1 net668 _10923__668/LO sky130_fd_sc_hd__conb_1
XFILLER_0_27_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06853__B2 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07163_ _02059_ _02773_ _02775_ _02072_ _02815_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06524__B net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06114_ net173 net141 net190 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__a21oi_1
X_07094_ _02737_ _02738_ _02740_ _02747_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06045_ net1088 _01633_ _01641_ _01730_ _01734_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[4\]
+ sky130_fd_sc_hd__a2111oi_2
Xclkbuf_leaf_62_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09555__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_4
Xfanout214 net216 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_4
XANTENNA__06540__A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout225 _04582_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout392_A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout236 net240 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_4
Xfanout247 _04824_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_2
X_09804_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\] _04811_ _04818_
+ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__and3_1
Xfanout258 net262 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_4
Xfanout269 _04805_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
X_07996_ net452 net715 vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__xor2_1
XANTENNA__07581__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__a31o_1
X_06947_ net201 _02500_ _02509_ _02617_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout180_X net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] _04721_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06878_ _02548_ _02546_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_55_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08617_ _04045_ net458 _04044_ vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05829_ _00712_ _01516_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__nand2_1
X_09597_ _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__inv_2
XANTENNA__06258__Y _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10093__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08548_ net1147 _03961_ _04002_ vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_46_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10824__500 vssd1 vssd1 vccd1 vccd1 _10824__500/HI net500 sky130_fd_sc_hd__conb_1
XANTENNA__07097__A1 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08479_ _03926_ _03949_ _03950_ _03753_ _03751_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__o32a_1
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10510_ clknet_leaf_18_wb_clk_i _00378_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10441_ clknet_leaf_46_wb_clk_i _00325_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_135_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10372_ clknet_leaf_22_wb_clk_i net726 net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_32_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05782__C_N _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout93_X net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07546__A _02235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06450__A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[44\]
+ vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07021__B2 team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06375__A3 _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05066__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06609__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07088__A1 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10708_ clknet_leaf_71_wb_clk_i _00539_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06625__A _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10639_ clknet_leaf_45_wb_clk_i _00503_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09936__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10992__633 vssd1 vssd1 vccd1 vccd1 _10992__633/HI net633 sky130_fd_sc_hd__conb_1
XFILLER_0_80_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06360__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09001__A2 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07850_ _01094_ net161 vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06801_ _01590_ _01598_ _02470_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__and3_1
X_07781_ _03281_ _03283_ _03299_ _03301_ _03276_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__o221a_1
X_04993_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1 vssd1
+ vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
Xinput3 gpio_in[24] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_2
X_09520_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\] _01420_
+ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__nand2_1
X_06732_ _02369_ _02378_ _02384_ _02404_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__or4b_1
XFILLER_0_78_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06663_ _02293_ _02294_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__or2_1
X_09451_ net919 net208 _04596_ vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08402_ _00711_ _03876_ _03854_ _03718_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__a211oi_1
X_05614_ net446 net444 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09382_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ _04541_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__nand3_1
XFILLER_0_59_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06594_ net258 _02265_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ team_07_WB.instance_to_wrap.team_07.circlePixel _03671_ net485 _00727_ vssd1
+ vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__o211ai_2
X_05545_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout238_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08264_ _00663_ _03704_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05476_ net299 _01018_ _01182_ _01184_ _01188_ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06535__A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07215_ _01795_ _01901_ _02865_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08195_ net485 _03673_ net489 vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__a21o_1
XANTENNA__06254__B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout405_A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07146_ _02793_ _02797_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07077_ net95 net89 net86 vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06028_ net171 _01715_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05317__C _01014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ _03308_ _03441_ _03533_ _03496_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__o31a_1
X_09718_ net1176 _04756_ _04757_ _04759_ vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990_ net631 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_87_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10640__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09649_ _00761_ _04712_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08644__B _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06817__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05987__C _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10976__617 vssd1 vssd1 vccd1 vccd1 _10976__617/HI net617 sky130_fd_sc_hd__conb_1
XFILLER_0_123_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10424_ clknet_leaf_12_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[1\]
+ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06045__A2 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10355_ clknet_leaf_56_wb_clk_i _00295_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09519__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10286_ clknet_leaf_5_wb_clk_i _00278_ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_104_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05067__Y _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06339__B _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06058__C _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05330_ _01036_ _01041_ vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08046__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09470__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05261_ _00973_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
X_07000_ _02662_ _02663_ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05192_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00904_ vssd1 vssd1
+ vccd1 vccd1 _00905_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07233__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07233__B2 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08951_ net490 _04242_ vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07902_ net258 _03456_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__or2_1
X_08882_ _01966_ _04203_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07914__A _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ _03381_ _03387_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout188_A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _03311_ _03312_ _03318_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__nand3_2
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04976_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] vssd1
+ vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
X_09503_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[21\]
+ net270 _04627_ _04629_ net223 vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__a221o_1
X_06715_ _01804_ _02044_ _02013_ net258 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__and4b_1
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07695_ _02109_ net82 _02771_ _01637_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout355_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09434_ _04556_ _03593_ _00813_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__mux2_1
XANTENNA__05153__B team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06646_ _02316_ _02317_ _02318_ _02313_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09365_ _04533_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__inv_2
X_06577_ _02178_ _02249_ _02250_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout143_X net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08316_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\] _03744_ _03780_
+ _03709_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05528_ _01238_ _01240_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__or2_1
X_09296_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ _04481_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09461__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05459_ _01167_ _01168_ _01170_ _01171_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__or4_1
X_08247_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\] _00730_ _03724_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\] vssd1 vssd1 vccd1 vccd1
+ _03726_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08178_ _00703_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__nand2_2
XFILLER_0_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07224__A1 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07224__B2 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ _02277_ _02758_ _02782_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__a21o_1
XANTENNA__06712__B _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10140_ clknet_leaf_32_wb_clk_i team_07_WB.instance_to_wrap.team_07.recPLAYER.playerDetect
+ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10071_ clknet_leaf_35_wb_clk_i _00129_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07824__A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05538__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06735__B1 _01413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10973_ net614 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06159__B _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05998__B net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06175__A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06606__C _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07558__X _03117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10407_ clknet_leaf_12_wb_clk_i _00298_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_104_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10338_ clknet_leaf_34_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.activate_rand_delay_2
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10269_ clknet_leaf_74_wb_clk_i _00261_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07734__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05254__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__B1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06500_ _02139_ _02160_ _02166_ _02032_ _02159_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07480_ _01961_ _03038_ _03039_ _03040_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_17_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06431_ _02062_ _02076_ _02104_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07900__C net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ _04379_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__inv_2
X_06362_ net136 net129 _01935_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__and3_4
XFILLER_0_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05313_ _01008_ _01025_ vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__nor2_1
X_08101_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[1\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__mux4_1
XFILLER_0_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06293_ net441 _01968_ _01967_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a21oi_2
X_09081_ _04328_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08032_ _00706_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ net295 _03567_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05244_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] _00956_ vssd1 vssd1
+ vccd1 vccd1 _00957_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07909__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05175_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\]
+ _00883_ vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08954__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09983_ clknet_leaf_83_wb_clk_i _00088_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05148__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08934_ net432 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ net241 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08299__X _03777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__A2 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ _04194_ _04193_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\] vssd1
+ vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__mux2_1
X_07816_ _03370_ _03368_ _03369_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__or3b_1
X_08796_ _04151_ _04152_ net195 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_84_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07747_ _03299_ _03301_ _03286_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__nand3b_1
X_04959_ net1178 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout260_X net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07678_ _03119_ _03153_ _03235_ _02697_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09417_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\]
+ _04570_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__nor2_1
X_06629_ _02164_ _02301_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ net226 _04519_ _04521_ net408 net881 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09279_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05456__B1 _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07819__A _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06723__A _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10123_ clknet_leaf_29_wb_clk_i _00161_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10054_ clknet_leaf_29_wb_clk_i net756 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input33_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06708__B1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05345__Y _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08937__X _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10956_ net597 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07133__B1 _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10887_ net563 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
XFILLER_0_85_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold108 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sdi vssd1 vssd1
+ vccd1 vccd1 net778 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_117_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10787__SET_B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold119 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_dc vssd1 vssd1
+ vccd1 vccd1 net789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06352__B _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09944__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06980_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _02643_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] vssd1 vssd1
+ vccd1 vccd1 _02646_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05931_ net287 _01623_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__nand2_4
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08650_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04077_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__xnor2_1
X_05862_ _01548_ _01555_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07601_ _03070_ _03093_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__or2_1
X_08581_ _04016_ _04024_ _03996_ vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_87_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_05793_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\] vssd1 vssd1
+ vccd1 vccd1 _01487_ sky130_fd_sc_hd__a41o_1
XFILLER_0_135_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07532_ _03084_ _03086_ _03090_ _03075_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06808__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07463_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ net395 net296 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ _03032_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[25\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07675__A1 _03162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06478__A2 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05396__C_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06527__B _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09202_ _04372_ _04413_ _04414_ _04416_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__or4_1
XFILLER_0_91_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06414_ _01675_ _01708_ net203 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__o21a_2
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07394_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[4\]
+ _02987_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__or4b_1
XFILLER_0_8_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06345_ _00710_ net132 _01698_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout318_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09064_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__or4_1
X_06276_ net183 _01929_ _01948_ _01952_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__o211a_1
XANTENNA__06543__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08015_ net1034 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_left
+ sky130_fd_sc_hd__and2b_1
X_05227_ _00883_ net301 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_102_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout106_X net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06262__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05158_ _00867_ _00868_ _00869_ _00870_ vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__a22o_1
XANTENNA__07077__C net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05089_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__or2_1
X_09966_ clknet_leaf_90_wb_clk_i _00071_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_08917_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__xnor2_1
X_09897_ _01777_ _04885_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ net298 net295 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ _04184_ vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08779_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\] net411 net982
+ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10810_ clknet_leaf_78_wb_clk_i _00631_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10741_ clknet_leaf_67_wb_clk_i _00571_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07666__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07130__A3 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10672_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[4\]
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05429__B1 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07969__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07549__A _02838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06453__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05069__A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07197__A3 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05356__X _01069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ clknet_leaf_55_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[3\]
+ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10037_ _00057_ _00648_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05904__A1 _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10939_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sck vssd1 vssd1
+ vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08854__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09939__A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10841__517 vssd1 vssd1 vccd1 vccd1 _10841__517/HI net517 sky130_fd_sc_hd__conb_1
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06130_ _01677_ _01692_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__nor2_4
XFILLER_0_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06363__A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06061_ _00685_ _00828_ _00959_ _00961_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__or4_4
X_05012_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] _00649_
+ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__nand2_2
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09820_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\] _04825_ _04833_
+ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__and3_1
Xfanout407 net410 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_2
Xfanout418 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_col vssd1 vssd1
+ vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06810__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout429 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_2
X_09751_ net248 _04780_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__nor2_1
X_06963_ _02479_ _02553_ _02633_ _02603_ _02557_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__a311o_1
X_08702_ _01241_ _04112_ _04114_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__and3_1
X_05914_ _00716_ net127 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__xnor2_1
X_09682_ _04732_ _04733_ _04735_ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__nor3_1
X_06894_ _02476_ _02528_ net115 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__a21oi_1
X_08633_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__nand2_1
XANTENNA__07922__A _01067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05845_ _01526_ _01529_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\]
+ _01523_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08564_ net140 _03962_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05776_ _01461_ _01467_ _01469_ _01474_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__nor4_4
XANTENNA__06538__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07515_ _02108_ _02150_ _03073_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__o21a_1
XANTENNA__07648__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08495_ _03630_ _03961_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07446_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\] _03021_
+ _02984_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06320__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07377_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\] _02977_
+ _02974_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07369__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09116_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ _04347_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__a31o_1
X_06328_ _01985_ _01990_ _01999_ _02003_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09047_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ _04299_ net252 vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__o21ai_1
X_06259_ net160 net150 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__nand2_8
XFILLER_0_32_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold450 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\] vssd1 vssd1
+ vccd1 vccd1 net1120 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold461 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\] vssd1 vssd1 vccd1
+ vccd1 net1131 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold472 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] vssd1 vssd1 vccd1
+ vccd1 net1153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06387__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09949_ net464 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_70_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10031__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07639__A1 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06167__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10724_ clknet_leaf_60_wb_clk_i _00554_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10655_ clknet_leaf_2_wb_clk_i _00510_ net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06454__Y _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__B _03857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload17 clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_16
XFILLER_0_51_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06183__A net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10586_ clknet_leaf_40_wb_clk_i _00450_ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.ssdec_ss
+ sky130_fd_sc_hd__dfstp_1
Xclkload28 clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_24_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload39 clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__inv_8
XFILLER_0_134_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05630_ _01331_ _01342_ _01337_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__or3b_1
XFILLER_0_99_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06358__A _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05561_ _01257_ _01264_ _01262_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07300_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__a21oi_1
X_08280_ _03637_ _03641_ _03657_ _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__or4_1
X_05492_ net422 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07231_ _02033_ _02775_ _02872_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07162_ net104 _02277_ _02767_ net166 vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06113_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _00710_ _01436_
+ _01434_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\] vssd1
+ vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__a32o_1
X_07093_ _02152_ _02742_ _02746_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold44_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06044_ net156 net124 _01732_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__o21ai_4
XANTENNA__06380__X _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout204 _01662_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06540__B net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout215 net216 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout226 _04510_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_2
Xfanout237 net239 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_4
X_09803_ _04821_ _04822_ vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__and2_1
Xfanout248 _04765_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_2
X_07995_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__xor2_1
Xfanout259 net262 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_2
X_09734_ net1153 _04769_ _04770_ vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__a21bo_1
XANTENNA__05156__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06946_ net217 _02510_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_31_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09665_ net1101 _04722_ _04723_ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__a21o_1
XANTENNA__07869__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ net93 _02545_ _02547_ _02472_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout173_X net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08616_ _01929_ _01926_ _00964_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__mux2_1
X_05828_ _01509_ _01520_ _01507_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__o21ai_1
X_09596_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\]
+ _04672_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06541__A1 _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06268__A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06541__B2 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08547_ _03610_ _04001_ net140 vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__a21o_1
X_05759_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08478_ net468 net472 _03664_ _03899_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__o311a_1
XFILLER_0_37_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07429_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\]
+ _03008_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\] vssd1
+ vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10440_ clknet_leaf_45_wb_clk_i net843 net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10371_ clknet_leaf_22_wb_clk_i net685 net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07827__A _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold280 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold291 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[1\]
+ vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06450__B _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout86_X net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05347__A _01000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07562__A _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06609__C _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10707_ clknet_leaf_71_wb_clk_i _00538_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06625__B _02119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10638_ clknet_leaf_43_wb_clk_i _00502_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10569_ clknet_leaf_26_wb_clk_i _00437_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06599__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05809__X _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06360__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06800_ _02466_ _02470_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_127_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07780_ _03279_ _03334_ _03274_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__o21bai_1
X_04992_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel vssd1 vssd1
+ vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
XANTENNA__06771__A1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 gpio_in[25] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_2
XFILLER_0_127_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06771__B2 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06731_ _02386_ _02387_ _02392_ _02400_ _02403_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06359__Y _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09450_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[2\]
+ net272 _04595_ net290 net220 vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a221o_1
X_06662_ _01639_ _02259_ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10847__523 vssd1 vssd1 vccd1 vccd1 _10847__523/HI net523 sky130_fd_sc_hd__conb_1
X_08401_ _03834_ _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05613_ net445 net444 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__and2_1
X_09381_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ _04538_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__a31o_1
X_06593_ net258 _02021_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08332_ _03805_ _03808_ net485 vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__a21o_1
X_05544_ net420 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 _01257_ sky130_fd_sc_hd__or3_2
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08263_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\] _03741_
+ net488 vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05475_ _01185_ _01186_ _01187_ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__or3b_1
XFILLER_0_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06535__B net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07214_ _02134_ net81 _02741_ _02861_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08194_ net416 team_07_WB.instance_to_wrap.team_07.circlePixel _03672_ vssd1 vssd1
+ vccd1 vccd1 _03673_ sky130_fd_sc_hd__or3b_1
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07145_ _02797_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07076_ _02726_ _02729_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06027_ net171 _01716_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__or2_1
XANTENNA__07539__B1 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10934__584 vssd1 vssd1 vccd1 vccd1 _10934__584/HI net584 sky130_fd_sc_hd__conb_1
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ net132 _03304_ _03474_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ _00655_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] vssd1
+ vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06929_ _02588_ _02590_ _02598_ _02599_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_87_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09648_ _00655_ _04709_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07711__B1 _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09579_ _01793_ _03967_ _03976_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_26_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09464__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07321__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06445__B net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10423_ clknet_leaf_13_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[0\]
+ net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_33_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10354_ clknet_leaf_56_wb_clk_i _00294_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06461__A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10285_ clknet_leaf_5_wb_clk_i _00277_ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06505__A1 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06636__A _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05260_ _00971_ _00972_ vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__nand2_2
XFILLER_0_127_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05191_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[24\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[26\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[28\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[30\]
+ _00899_ _00900_ vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__mux4_2
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07233__A2 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06371__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08950_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _00710_ _04234_
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_cleared vssd1 vssd1 vccd1 vccd1
+ _04242_ sky130_fd_sc_hd__a31o_1
X_07901_ _01058_ net216 _01723_ _03384_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__o22a_1
X_08881_ net1081 _04205_ vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07832_ _03382_ _03385_ _03386_ _03375_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__or4b_2
XFILLER_0_138_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07763_ _03317_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__inv_2
X_10888__645 vssd1 vssd1 vccd1 vccd1 net645 _10888__645/LO sky130_fd_sc_hd__conb_1
X_04975_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\] vssd1
+ vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
X_09502_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\] vssd1
+ vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06714_ _02135_ _02259_ _02312_ _02140_ _02221_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07694_ net111 _03249_ _01639_ _02760_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__or4b_1
XFILLER_0_91_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09433_ _04557_ _03592_ _00813_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__mux2_2
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06645_ net286 _00757_ _02297_ _02308_ _02109_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout348_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09364_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ _04530_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06576_ net93 net108 net95 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_74_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08315_ _03695_ _03792_ _03738_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a21oi_1
X_05527_ _01239_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__nand2b_2
X_09295_ net229 _04483_ _04484_ net404 net1068 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__a32o_1
XANTENNA_20 _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_31 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout136_X net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08246_ _01284_ _01305_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__nand2_1
X_05458_ _01002_ _01016_ _01035_ _01099_ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__or4_1
XANTENNA__07472__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08177_ net471 _03655_ net469 vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05389_ _00966_ _00967_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07128_ _02761_ _02764_ _02768_ _02781_ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07224__A2 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06712__C _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07059_ _01630_ _02212_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10070_ clknet_leaf_35_wb_clk_i _00128_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07543__C net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10424__RESET_B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06684__A_N _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10972_ net613 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
XANTENNA__08488__B2 net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06175__B net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10406_ clknet_leaf_11_wb_clk_i net716 net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08412__A1 _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10337_ clknet_leaf_51_wb_clk_i net676 net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_108_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10268_ clknet_leaf_74_wb_clk_i _00260_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07734__B _01104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ clknet_leaf_86_wb_clk_i _00203_ net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06726__A1 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05934__C1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10165__RESET_B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05254__B team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07750__A _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05822__X _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07151__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07151__B2 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06430_ _02092_ _02103_ _02090_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08057__S net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06366__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06361_ net163 _01653_ _01685_ _01683_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08100_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[4\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[5\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[6\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[7\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__mux4_1
X_05312_ _00996_ _01010_ vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__or2_2
XFILLER_0_86_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06292_ net438 net440 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08031_ net455 net452 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05243_ _00953_ _00954_ _00955_ _00947_ vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__o31a_1
Xinput40 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05174_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00886_ vssd1 vssd1
+ vccd1 vccd1 _00887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06414__B1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08954__A2 _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09982_ clknet_leaf_83_wb_clk_i _00087_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[17\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07484__X _03045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06965__B2 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08933_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] net1142 net242 vssd1
+ vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__mux2_1
XANTENNA__06666__A2_N _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout298_A _03026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08864_ net450 net263 _04192_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__and3_1
X_07815_ _01057_ _01741_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__nor2_1
X_08795_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\] _04147_ net959
+ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout465_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07746_ _03290_ _03300_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__and2_1
X_04958_ net1134 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ net202 _01723_ _01736_ _02829_ _03217_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout253_X net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ _04568_ _04569_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06628_ _02296_ _02300_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09347_ _04520_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06559_ _02228_ _02230_ _02232_ _02227_ _02226_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ _04264_ net228 _04472_ net401 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__a32o_1
XANTENNA__08491__A net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06653__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08229_ net416 _03707_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07819__B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10122_ clknet_leaf_28_wb_clk_i _00160_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07835__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ clknet_leaf_30_wb_clk_i net772 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06708__B2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05355__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10955_ net596 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_74_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10886_ net562 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_39_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold109 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06947__A1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05930_ net286 net278 _01621_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07464__B net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05861_ _01538_ _01554_ _01542_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__mux2_2
X_07600_ _03069_ _03097_ _03125_ _03158_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_1_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08580_ _03619_ _04023_ net139 vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05792_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__nand4_4
XFILLER_0_44_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07480__A _01961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07531_ _03081_ _03087_ _03089_ _02034_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__and4b_1
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07124__B2 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06808__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07462_ net454 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09201_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__or4_1
X_06413_ net137 net105 net169 _02086_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a31o_2
XANTENNA__06527__C _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07393_ _02988_ _02989_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_33_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09132_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ _04327_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__or3_1
X_06344_ net418 net134 _02016_ _02018_ net128 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09063_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__or4b_1
XFILLER_0_5_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06275_ _01931_ _01949_ _01950_ _01951_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08014_ net1007 net729 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_down
+ sky130_fd_sc_hd__and2b_1
X_05226_ _00685_ _00938_ _00828_ _00928_ vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__or4b_1
XFILLER_0_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08927__A2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05157_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00870_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05088_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__nor2_2
X_09965_ clknet_leaf_87_wb_clk_i _00070_ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_110_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08916_ _00724_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_x\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[2\]
+ _00725_ _04224_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__a221o_1
X_09896_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[9\] _01776_ vssd1
+ vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ net396 net394 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\]
+ net411 vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__or3_1
XANTENNA__06558__X _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05462__X _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05903__A _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07729_ _03277_ _03283_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07115__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10740_ clknet_leaf_72_wb_clk_i _00570_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07666__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08863__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[3\]
+ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05069__B _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10105_ clknet_leaf_55_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[2\]
+ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09879__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10036_ _00056_ _00647_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10141__D team_07_WB.instance_to_wrap.team_07.recFLAG.flagDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05904__A2 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10938_ team_07_WB.instance_to_wrap.ssdec_sck vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10869_ net545 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_27_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10880__556 vssd1 vssd1 vccd1 vccd1 _10880__556/HI net556 sky130_fd_sc_hd__conb_1
XFILLER_0_54_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06363__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06060_ _01457_ _01481_ _01483_ _00653_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_1_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05011_ _00635_ net288 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout408 net410 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_2
Xfanout419 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[11\] vssd1
+ vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_2
XANTENNA__08790__B1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10180__RESET_B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ _04767_ _04780_ _04781_ net249 net1131 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__a32o_1
X_06962_ _02483_ _02632_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__nand2_1
X_08701_ _04120_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ _04115_ vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__mux2_1
X_05913_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] net127
+ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__xnor2_2
X_09681_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ net250 vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__and3_1
X_06893_ net111 _02563_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07345__B2 _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04059_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__nand2_1
XANTENNA__07922__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05844_ _01534_ _01537_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08563_ _03614_ _04011_ net139 vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__a21oi_1
X_05775_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\]
+ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout163_A _01557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07514_ net100 _02191_ _03072_ _01612_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ _03962_ net53 _03961_ vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__mux2_1
XANTENNA__07648__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07445_ _03021_ _03022_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[22\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout330_A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07376_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\] _02977_
+ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09115_ net212 _04352_ _04353_ net400 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06327_ _01987_ _01989_ _02002_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06273__B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout216_X net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09046_ _00664_ _04300_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06258_ net157 net145 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__nor2_2
XFILLER_0_128_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05209_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00922_ sky130_fd_sc_hd__nand2_1
Xhold440 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[0\] vssd1 vssd1
+ vccd1 vccd1 net1110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06189_ net289 net134 _01848_ _01861_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a211o_1
Xhold451 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold473 team_07_WB.instance_to_wrap.team_07.label_num_bus\[28\] vssd1 vssd1 vccd1
+ vccd1 net1143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[21\]
+ vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06387__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07584__A1 _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09948_ net464 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_70_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09879_ net837 net153 net151 _04874_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07324__S _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08647__C _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06448__B _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10723_ clknet_leaf_60_wb_clk_i _00553_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06847__B1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10654_ clknet_leaf_2_wb_clk_i _00509_ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_24_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06464__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08064__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10585_ clknet_leaf_53_wb_clk_i _00449_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload18 clknet_leaf_81_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__inv_12
XANTENNA__06183__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload29 clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_23_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_114_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08772__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ clknet_leaf_42_wb_clk_i _00098_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_99_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05560_ _01270_ _01271_ _01269_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__o21bai_1
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05491_ _01198_ _01200_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07230_ net129 net141 _02773_ _02877_ _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__a41o_1
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10779__RESET_B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07161_ _02793_ _02798_ _02811_ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06112_ _00827_ _01789_ _01794_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__a22o_1
XANTENNA__06524__D _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07092_ _01654_ net164 _01664_ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06043_ net156 net124 _01732_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05718__A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 _01661_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_4
Xfanout216 _01503_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_4
Xfanout227 _04510_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_2
X_09802_ _04811_ _04818_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__a21o_1
Xfanout238 net239 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_4
Xfanout249 _04765_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_1
X_07994_ _03546_ _03547_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__xnor2_1
X_09733_ _00652_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[2\] net248
+ _04768_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__or4_1
X_06945_ net257 _02508_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__nor2_1
X_09664_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] _04719_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\] vssd1 vssd1 vccd1
+ vccd1 _04723_ sky130_fd_sc_hd__and4b_1
X_06876_ _01590_ _01598_ _02470_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07869__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08615_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] _04044_ vssd1 vssd1
+ vccd1 vccd1 _00176_ sky130_fd_sc_hd__xnor2_1
X_05827_ _01513_ _01516_ _00712_ _01507_ _01509_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__a2111o_1
X_09595_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\] _04672_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_71_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout166_X net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08546_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ _03608_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__o21ai_1
X_05758_ _01454_ _01455_ _01456_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_46_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08477_ _03898_ _03948_ _03667_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__o21a_1
X_05689_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[0\] team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[1\]
+ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[2\] team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[3\]
+ net441 net440 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07428_ net966 _03009_ _03011_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[16\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_98_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06284__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06715__C _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07359_ net1180 _02965_ _02967_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__or4b_1
XFILLER_0_61_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10904__570 vssd1 vssd1 vccd1 vccd1 _10904__570/HI net570 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_135_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10370_ clknet_leaf_23_wb_clk_i net699 net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09029_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ _04286_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07827__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[11\] vssd1 vssd1
+ vccd1 vccd1 net940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09546__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold281 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] vssd1 vssd1
+ vccd1 vccd1 net951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08939__A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05915__X _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06780__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05363__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10706_ clknet_leaf_70_wb_clk_i _00537_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10637_ clknet_leaf_43_wb_clk_i _00501_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10568_ clknet_leaf_27_wb_clk_i _00436_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06599__A2 _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10499_ clknet_leaf_16_wb_clk_i _00367_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06641__B _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05257__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07753__A _01067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04991_ team_07_WB.instance_to_wrap.team_07.lcdOutput.stagePixel vssd1 vssd1 vccd1
+ vccd1 _00728_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput5 gpio_in[26] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06730_ _02402_ _02397_ _02394_ _02401_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_36_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06661_ _02108_ _02259_ _02333_ net89 net98 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__o221a_1
X_10886__562 vssd1 vssd1 vccd1 vccd1 _10886__562/HI net562 sky130_fd_sc_hd__conb_1
X_08400_ _03738_ _03871_ _03874_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__o21a_1
X_05612_ net446 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__and2b_1
X_09380_ net226 _04543_ _04544_ net409 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__a32o_1
X_06592_ _02021_ _01654_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08331_ _00729_ _03736_ _03807_ _03738_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05543_ net420 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 _01256_ sky130_fd_sc_hd__nor3_2
XFILLER_0_15_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08262_ _00728_ _03740_ _03700_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__a21o_1
X_05474_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ net192 _01021_ _01062_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07213_ _02073_ _02862_ _02863_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08193_ team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel team_07_WB.instance_to_wrap.team_07.borderGen.borderPixel
+ team_07_WB.instance_to_wrap.team_07.flagPixel vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout126_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07144_ _02794_ _02796_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07075_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\] net301 net300 team_07_WB.instance_to_wrap.team_07.label_num_bus\[24\]
+ _02728_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a221o_2
X_06026_ net171 _01716_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__nor2_1
XANTENNA__07539__A1 _02080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _00747_ _03414_ _03416_ _00746_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__o22a_1
X_09716_ _04757_ _04758_ vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__and2_1
X_06928_ net133 _02497_ _02503_ _02596_ _02521_ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a41o_1
XFILLER_0_97_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ _04703_ _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06859_ net115 _02471_ _02529_ net108 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__o22a_1
XANTENNA__07711__A1 _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06514__A2 _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _04637_ _04661_ net480 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ net1005 _03988_ vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_137_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06445__C net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10422_ clknet_leaf_13_wb_clk_i net242 net334 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07838__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10353_ clknet_leaf_59_wb_clk_i _00293_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06461__B _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ clknet_leaf_5_wb_clk_i _00276_ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.stage\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06202__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913__658 vssd1 vssd1 vccd1 vccd1 net658 _10913__658/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_109_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07702__A1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06269__A1 _00684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06269__B2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07748__A _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05190_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00901_ vssd1 vssd1
+ vccd1 vccd1 _00903_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07610__A2_N _03144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08718__B1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07900_ _03384_ _03454_ net256 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__and3b_1
XFILLER_0_110_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08880_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_cleared _04204_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__or3b_1
X_07831_ _01094_ net186 vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__nor2_1
X_07762_ _01076_ net189 _03316_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__a21o_1
X_04974_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\] vssd1
+ vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09501_ net926 net206 _04628_ vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__o21a_1
X_06713_ _01732_ _02283_ _02385_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__o21a_1
X_07693_ _00759_ net119 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__and2_1
XANTENNA__09694__A1 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10410__Q team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09432_ net1155 _04578_ _04579_ _04581_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__o22a_1
X_06644_ _02164_ _02295_ _02301_ _01921_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09363_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ _04530_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__or2_1
X_06575_ _00754_ _02138_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout243_A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07457__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05526_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ _01196_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__and2_1
X_08314_ _03791_ _01302_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__mux2_1
X_09294_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ _04481_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__or2_1
XANTENNA_10 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_21 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_32 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08245_ _01285_ _01306_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05457_ net435 _01072_ _01113_ _01036_ _01169_ vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout410_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout129_X net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08176_ net474 net472 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__nor2_1
XANTENNA__06562__A _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05388_ _01099_ _01100_ _01066_ vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07127_ _00755_ net86 _02780_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__a21oi_4
XANTENNA__07224__A3 _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07058_ _01630_ _02209_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__nor2_1
XANTENNA__06712__D _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06009_ net134 net143 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08489__A net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input3_X net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10971_ net612 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_69_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10982__623 vssd1 vssd1 vccd1 vccd1 _10982__623/HI net623 sky130_fd_sc_hd__conb_1
XANTENNA__05912__Y _01606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07840__B net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07332__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07568__A _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10405_ clknet_leaf_10_wb_clk_i net689 net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_68_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10336_ clknet_leaf_51_wb_clk_i net672 net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10267_ clknet_leaf_74_wb_clk_i _00259_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10198_ clknet_leaf_83_wb_clk_i _00202_ net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06726__A2 _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05934__B1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07750__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06647__A _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07151__A2 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06366__B _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06360_ net131 net126 _01686_ _01936_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__or4_2
XFILLER_0_17_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05311_ net191 _01015_ _01023_ vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_86_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06291_ net438 _01397_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08030_ _03566_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net393 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__mux2_1
X_05242_ net301 _00874_ _00900_ net300 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__a22o_1
XANTENNA__07478__A _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput30 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput41 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06382__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05173_ _00884_ _00885_ _00873_ vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06414__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07611__B1 _01672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09981_ clknet_leaf_83_wb_clk_i _00086_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_12_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08932_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ net241 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08167__A1 net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08863_ net450 _04192_ _04193_ vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07814_ _01113_ net186 vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__nand2_1
X_08794_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\]
+ _04147_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__or3_1
X_10966__607 vssd1 vssd1 vccd1 vccd1 _10966__607/HI net607 sky130_fd_sc_hd__conb_1
XANTENNA__07941__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04957_ net7 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07745_ _00753_ _03292_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout360_A net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout458_A team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07676_ _02040_ _02260_ _03198_ _01655_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09415_ net481 _02961_ _04556_ _00819_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10305__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06627_ _02265_ _02294_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout246_X net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09346_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ _04514_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__and3_1
X_06558_ net121 net204 _02231_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05509_ net424 net423 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__and2b_1
X_09277_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06489_ _02155_ _02162_ _02161_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08228_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03706_ vssd1
+ vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08159_ net475 _03640_ _03642_ _03638_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05339__C _01005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10121_ clknet_leaf_28_wb_clk_i _00159_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07327__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ clknet_leaf_29_wb_clk_i net787 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05355__B _01067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07851__A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input19_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10954_ net595 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_98_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07133__A2 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10885_ net561 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_35_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06892__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06644__A1 _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06644__B2 _01921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09594__B1 _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10919__664 vssd1 vssd1 vccd1 vccd1 net664 _10919__664/LO sky130_fd_sc_hd__conb_1
XFILLER_0_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ clknet_leaf_47_wb_clk_i net744 net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__05546__A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05860_ _01534_ _01536_ _01537_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05791_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] vssd1 vssd1
+ vccd1 vccd1 _01485_ sky130_fd_sc_hd__nand3_1
XANTENNA__06580__B1 _02230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07530_ net181 net171 _02082_ _02097_ _03088_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__o311a_1
XFILLER_0_44_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07461_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ net396 net297 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ _03031_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[24\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06332__B1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09200_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__or4b_1
X_06412_ net214 net138 _01706_ _02054_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a31oi_4
X_07392_ net1177 _02987_ net480 vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06343_ _01724_ _02012_ _02017_ _02011_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__or4b_1
X_09131_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ _04318_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__nand3_1
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06824__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09062_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__or2_1
XANTENNA__05438__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06274_ _00684_ net458 net201 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05225_ _00935_ _00936_ _00937_ _00931_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__o31a_1
X_08013_ net1001 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_up
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout206_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05156_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07936__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07060__A1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05087_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[2\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[1\]
+ _00812_ vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__or3_2
X_09964_ clknet_leaf_88_wb_clk_i _00069_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_34_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09337__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__xor2_1
X_09895_ net844 net154 net152 _04884_ vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout196_X net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ net749 _04183_ vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__and2_1
XANTENNA__06804__A1_N net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08777_ _04138_ net411 net1105 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__mux2_1
X_05989_ _01677_ _01679_ net171 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05903__B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07728_ _01065_ net120 vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__nor2_1
XANTENNA__07115__A2 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07659_ _01680_ net167 _02835_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07666__A3 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10670_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[2\]
+ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09329_ _00662_ _04507_ _04508_ _04503_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08076__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06626__A1 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09576__B1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07051__A1 _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10104_ clknet_leaf_55_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[1\]
+ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_10035_ _00055_ _00646_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_19_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06909__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10937_ team_07_WB.instance_to_wrap.ssdec_ss vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10868_ net544 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_73_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08616__S _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10770__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10799_ clknet_leaf_73_wb_clk_i _00620_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06617__A1 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05010_ team_07_WB.EN_VAL_REG net41 _00745_ vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__mux2_1
XANTENNA__06660__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout409 net410 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_120_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06961_ _00695_ _02106_ _00749_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08700_ _04117_ _04118_ _04119_ net263 vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__o211a_1
X_05912_ _01596_ _01603_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09680_ _00655_ _04703_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nand2_1
XANTENNA__06659__X _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06892_ net434 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] _02466_ _02467_
+ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__o22a_1
X_08631_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__or3b_2
X_05843_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] _01520_
+ _01523_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__and3_1
X_08562_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[10\]
+ _03613_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__o21ai_1
X_05774_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[11\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\] _01472_ vssd1
+ vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__or4b_1
XANTENNA__06160__A1_N net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07513_ net94 _01629_ _02332_ net96 vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__a31o_1
X_08493_ _03650_ _03652_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout156_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07444_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\] _03019_
+ net478 vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07375_ _02977_ _02978_ _02974_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[3\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout323_A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09114_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ _04350_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06326_ net218 _01969_ _02000_ _02001_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09045_ net252 _04298_ _04300_ net403 net1066 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06257_ _01933_ _01925_ _01923_ _01932_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__nand4b_1
XTAP_TAPCELL_ROW_96_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout111_X net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout209_X net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05208_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00921_ sky130_fd_sc_hd__or2_1
Xhold430 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06188_ _01852_ _01868_ _01854_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a21oi_1
Xhold441 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\] vssd1 vssd1
+ vccd1 vccd1 net1111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07033__A1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[2\] vssd1 vssd1
+ vccd1 vccd1 net1133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05139_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00852_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\] vssd1 vssd1
+ vccd1 vccd1 net1144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold496 team_07_WB.instance_to_wrap.team_07.label_num_bus\[9\] vssd1 vssd1 vccd1
+ vccd1 net1166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06387__A3 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09947_ net464 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09878_ _01772_ _04873_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08829_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] _04141_
+ net1099 vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10722_ clknet_leaf_67_wb_clk_i _00010_ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05920__Y _01614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08049__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10653_ clknet_leaf_2_wb_clk_i _00508_ net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06464__B net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10584_ clknet_leaf_52_wb_clk_i _00448_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_24_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload19 clknet_leaf_83_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__inv_8
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09549__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06480__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07024__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10660__RESET_B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06479__X _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ clknet_leaf_42_wb_clk_i _00097_ net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[9\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10369__SET_B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05490_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ _01202_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07160_ _02058_ _02120_ _02812_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06111_ _01789_ _01793_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07091_ net255 _01657_ _01667_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06042_ net161 _01653_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__nand2_8
XFILLER_0_50_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout206 net209 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
X_09801_ _04811_ _04820_ _04808_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__a21o_1
Xfanout217 _01503_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05467__A_N _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout228 _04471_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
X_07993_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__xor2_1
X_09732_ net1151 _04766_ _04769_ vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06944_ net182 _02612_ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09663_ net1061 _04720_ _04722_ vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__o21a_1
XANTENNA__06526__B1 _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ net90 _02544_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout273_A _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ _04042_ _04043_ _00960_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__a21o_1
X_05826_ _01513_ _01516_ _00712_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__a21o_1
X_09594_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\] _04664_ _04666_
+ _04673_ vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08545_ _03609_ _04000_ _03999_ vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__a21oi_1
X_05757_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[18\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] _01453_ vssd1 vssd1
+ vccd1 vccd1 _01456_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout159_X net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ _03755_ _03819_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05688_ _00681_ net440 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07427_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\] _03009_
+ net233 vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_40_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_63_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06715__D net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07358_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\]
+ _02966_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_135_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08780__A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06057__A2 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06309_ net173 _01973_ _01984_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07289_ net442 _01326_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09028_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ _04286_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold260 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[2\]
+ vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10418__RESET_B net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[1\] vssd1
+ vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10831__507 vssd1 vssd1 vccd1 vccd1 _10831__507/HI net507 sky130_fd_sc_hd__conb_1
XANTENNA__07335__S _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950__591 vssd1 vssd1 vccd1 vccd1 _10950__591/HI net591 sky130_fd_sc_hd__conb_1
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06475__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10705_ clknet_leaf_68_wb_clk_i _00536_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07493__A1 _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10636_ clknet_leaf_44_wb_clk_i net880 net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10567_ clknet_leaf_26_wb_clk_i _00435_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10498_ clknet_leaf_16_wb_clk_i _00366_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10159__RESET_B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06360__D _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07753__B _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04990_ net416 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
Xinput6 gpio_in[27] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_3_4_0_wb_clk_i_X clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06660_ net283 net88 _02031_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05611_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\] net443
+ net444 _01323_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__o32a_1
XFILLER_0_8_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06591_ net123 _01654_ _02261_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__or3_2
XANTENNA__05731__A1 _00709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08330_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\] _03734_ _03806_
+ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05542_ net419 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] vssd1 vssd1 vccd1
+ vccd1 _01255_ sky130_fd_sc_hd__or3_2
XANTENNA__06385__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07484__A1 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08261_ team_07_WB.instance_to_wrap.team_07.buttonPixel team_07_WB.instance_to_wrap.team_07.buttonHighlightPixel
+ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__nor2_1
X_05473_ _01036_ _01037_ _01106_ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07212_ _01653_ _01665_ net188 vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_41_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08192_ team_07_WB.instance_to_wrap.team_07.flagPixel team_07_WB.instance_to_wrap.team_07.lcdOutput.playerPixel
+ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_41_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07143_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] net302 net398 _02795_
+ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06391__Y _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout119_A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[32\] net302 net398 _02727_
+ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a22o_1
XANTENNA__05729__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06025_ net218 net197 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07539__A2 _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _03280_ _03522_ _03530_ _03515_ _03518_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__o2111a_1
X_09715_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] net250 _04752_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\] vssd1 vssd1 vccd1
+ vccd1 _04758_ sky130_fd_sc_hd__a31o_1
X_06927_ _02593_ _02594_ _02596_ _02597_ _02589_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout276_X net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09646_ _01767_ _04709_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06858_ net434 _02528_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05809_ _01494_ _01499_ _01500_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__or3_4
X_09577_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\] _04661_
+ _04663_ _04640_ vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_26_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ _02410_ _02415_ _02460_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_26_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08528_ net1114 _03987_ vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_137_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06295__A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08459_ _03714_ _03749_ _03751_ _03931_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08941__C _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07227__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ clknet_leaf_56_wb_clk_i _00312_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07227__B2 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10352_ clknet_leaf_56_wb_clk_i _00292_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05789__B2 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05358__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10283_ clknet_leaf_86_wb_clk_i _00275_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07163__B1 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06476__Y _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09455__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06269__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07218__A1 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10619_ clknet_leaf_48_wb_clk_i _00483_ net373 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07748__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07830_ _03383_ _03384_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__or2_1
X_07761_ _03314_ _03315_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__nand2b_1
X_04973_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[10\] vssd1
+ vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
X_09500_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[20\]
+ net270 _04625_ _04627_ net220 vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a221o_1
X_06712_ net254 _01734_ _02021_ _02154_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07692_ _03041_ _03247_ _03248_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recMOD.modSquaresDetect
+ sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09431_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ _04569_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__and2b_1
X_06643_ _02031_ _02281_ _02314_ _02315_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__o211ai_1
XANTENNA__06386__Y _02060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09362_ net227 _04529_ _04531_ net409 net1063 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06574_ _02075_ _02098_ _02247_ net253 net87 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__o311a_1
XFILLER_0_87_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08313_ _01381_ _03733_ _03789_ _03790_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a2bb2o_1
X_05525_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ _01237_ _01236_ _01234_ _01194_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__a2111oi_4
X_09293_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ _04481_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__nand2_1
XANTENNA_11 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07498__X _03058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08244_ net485 net416 _03721_ net489 vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__a211o_1
XANTENNA_33 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[5\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05456_ _01006_ _01056_ _01063_ _01058_ _01052_ vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06843__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08175_ _00733_ net130 vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__nor2_1
X_05387_ net191 _01014_ _01021_ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout403_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06562__B _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08957__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07126_ net284 _00749_ net120 _01634_ _02779_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__a311o_1
XFILLER_0_43_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07057_ _01811_ _02036_ _02709_ _02711_ _01903_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06008_ net131 _01698_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__nor2_2
XANTENNA__05786__A4 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07959_ _00970_ _01058_ net117 _03513_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__a31o_1
XANTENNA__05943__A1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10970_ net611 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09629_ net1003 _04696_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__xor2_1
XANTENNA__06499__A2 _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06737__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05360__C _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08951__A_N net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06120__A1 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10048__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.idle vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07568__B _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10433__RESET_B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08948__A1 _00709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10404_ clknet_leaf_10_wb_clk_i net680 net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10335_ clknet_leaf_51_wb_clk_i net674 net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10837__513 vssd1 vssd1 vccd1 vccd1 _10837__513/HI net513 sky130_fd_sc_hd__conb_1
X_10266_ clknet_leaf_74_wb_clk_i _00258_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10197_ clknet_leaf_90_wb_clk_i _00201_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06726__A3 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05934__A1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07151__A3 _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05310_ _01003_ _01010_ _01021_ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__nor3_2
XFILLER_0_71_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06290_ _01397_ _01399_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__nand2_2
XFILLER_0_127_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05241_ net449 _00843_ net398 _00832_ vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__a31o_1
Xinput20 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput31 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05172_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\]
+ _00883_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10894__651 vssd1 vssd1 vccd1 vccd1 net651 _10894__651/LO sky130_fd_sc_hd__conb_1
XFILLER_0_12_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06414__A2 _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07611__A1 _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09980_ clknet_leaf_87_wb_clk_i _00085_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_122_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08931_ net434 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[0\]
+ net242 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08862_ net450 net240 _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__o21ai_1
XANTENNA__05726__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ _01112_ net189 _01658_ _01057_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__a22o_1
X_08793_ _04149_ _04150_ net196 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout186_A _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07744_ _01064_ net109 _03280_ _03284_ _01609_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_84_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04956_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1 vssd1 vccd1
+ vccd1 _00696_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07675_ _03162_ _03226_ _03232_ _03076_ _03225_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__a221o_1
XANTENNA__07678__B2 _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout353_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09414_ net477 _02961_ _04557_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06626_ _02109_ _02295_ _02297_ _02298_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a22oi_2
X_09345_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ _04514_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06557_ _01654_ _01829_ net205 vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout141_X net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_X net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07669__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05508_ _00691_ _01198_ _01203_ _00692_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__a22o_1
X_09276_ net228 net401 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06488_ _01655_ _02056_ _02054_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__o21a_1
XFILLER_0_106_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08227_ net2 _03704_ _03705_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__a31o_2
XFILLER_0_16_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05439_ _01151_ _01126_ _00965_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08158_ _03640_ _03642_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07109_ _01694_ net164 _02758_ _02761_ _02762_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08089_ _03597_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[9\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10120_ clknet_leaf_27_wb_clk_i _00158_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05917__A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout99_A _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10051_ clknet_leaf_29_wb_clk_i _00109_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06748__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10953_ net594 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_74_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10884_ net560 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06892__A2 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07624__A2_N _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08397__A2 _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07585__Y _03144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10318_ clknet_leaf_54_wb_clk_i net777 net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10249_ clknet_leaf_82_wb_clk_i _00241_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07109__B1 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05790_ net1037 _00797_ _00827_ net476 vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a22o_1
XANTENNA__06580__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07480__C _03039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07460_ net455 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06411_ net138 _01691_ net168 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__and3_2
XFILLER_0_57_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10355__RESET_B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07391_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[3\] _02987_
+ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09130_ net403 _04324_ _04363_ vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_33_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06342_ _00710_ net218 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__04906__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ _04309_ _04311_ _04307_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06273_ net458 net217 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08012_ _03558_ _03559_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__xnor2_1
X_05224_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00937_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09034__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05155_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00868_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout101_A _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05086_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[7\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[5\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[8\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__or4_1
X_09963_ clknet_leaf_84_wb_clk_i _00068_ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_65_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08914_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__xor2_1
X_09894_ _01776_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07952__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08845_ _04182_ _04183_ _04144_ vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_51_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06020__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_X net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ net411 _01457_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__nor2_1
XANTENNA__06571__A1 _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05988_ net189 net179 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__or2_2
X_07727_ _01064_ net116 _03281_ _03276_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__o31a_1
XFILLER_0_68_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_04939_ net442 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06287__B net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07658_ _01902_ _02087_ _03213_ _03215_ _03119_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__a32o_1
XFILLER_0_95_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06609_ net161 net127 _01652_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__and3_2
XFILLER_0_76_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10096__RESET_B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07589_ net255 _03146_ _03147_ _03145_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09328_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[16\]
+ net402 _04259_ net228 vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__a22o_1
XANTENNA__09273__A0 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06087__B1 _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09259_ _04458_ _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07338__S team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07051__A2 _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10103_ clknet_leaf_55_wb_clk_i team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[0\]
+ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_8_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input31_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _00054_ _00645_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_19_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10936_ team_07_WB.instance_to_wrap.ssdec_sdi vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10867_ net543 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05716__A_N net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10798_ clknet_leaf_78_wb_clk_i _00619_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07102__A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06363__D _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06660__B net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05557__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06005__X _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06960_ _02602_ _02604_ _02630_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05911_ _01597_ _01604_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__nand2_1
X_06891_ _02556_ _02561_ _02543_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a21o_1
XANTENNA__08587__B net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08630_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04046_ _04057_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05842_ _01527_ _01535_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__and2_1
XANTENNA__06388__A _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05292__A _00675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08561_ net140 _04010_ _03963_ vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__o21ai_1
X_05773_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[10\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__and4b_1
X_07512_ _01628_ _03070_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__or2_1
X_08492_ net1147 _03961_ vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06675__X _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload88_A clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07443_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\]
+ _03018_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout149_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07374_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__a31o_1
XANTENNA__09211__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09113_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ _04350_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__or2_1
X_06325_ net261 _01397_ net439 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__or3b_1
XFILLER_0_95_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout316_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09044_ _04299_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__inv_2
X_06256_ _00684_ net180 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_96_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05207_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00920_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold420 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\] vssd1 vssd1
+ vccd1 vccd1 net1090 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout104_X net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold431 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] vssd1 vssd1
+ vccd1 vccd1 net1101 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ _01855_ _01867_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold442 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold453 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[10\] vssd1 vssd1
+ vccd1 vccd1 net1134 sky130_fd_sc_hd__dlygate4sd3_1
X_05138_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00851_ sky130_fd_sc_hd__or2_1
XANTENNA__07033__A2 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold475 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[3\] vssd1 vssd1 vccd1
+ vccd1 net1156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09946_ net463 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
X_05069_ net492 _00796_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06792__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[2\] vssd1 vssd1 vccd1
+ vccd1 _04873_ sky130_fd_sc_hd__o21ai_1
X_08828_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\]
+ _04141_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__or3_1
XANTENNA__05914__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06544__A1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06298__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08759_ net902 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ net235 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05930__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10721_ clknet_leaf_62_wb_clk_i _00552_ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08049__A1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10652_ clknet_leaf_2_wb_clk_i _00507_ net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09246__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ clknet_leaf_53_wb_clk_i _00447_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10318__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06480__B net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07592__A _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ clknet_leaf_42_wb_clk_i _00096_ net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[8\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05824__B _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06001__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10919_ net664 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_128_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06110_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[8\] _01792_ vssd1 vssd1
+ vccd1 vccd1 _01793_ sky130_fd_sc_hd__and4b_2
XFILLER_0_41_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07090_ net255 _01657_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__nand2_4
XANTENNA__08460__A1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06671__A _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06041_ net158 _01652_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05287__A _00675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09800_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[5\] _04818_ vssd1
+ vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__nand2_1
Xfanout207 net209 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__buf_2
Xfanout218 net219 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_8
Xfanout229 _04471_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_2
X_07992_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ net1161 vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09731_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _04768_ net248
+ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a21o_1
X_06943_ net182 _02612_ _02613_ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10717__RESET_B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09662_ _04716_ _04721_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__nor2_1
X_06874_ _02544_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__inv_2
XANTENNA__07723__B1 _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ _00964_ _01927_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__nand2_1
X_05825_ _00712_ net200 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__nor2_1
XANTENNA__10370__RESET_B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09593_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\] _04672_ vssd1
+ vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08544_ net862 _03608_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__nand2_1
X_05756_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[21\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[20\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\] vssd1 vssd1 vccd1
+ vccd1 _01455_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08475_ _03908_ _03946_ net491 _03753_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_46_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05687_ _00681_ net440 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07426_ _03009_ _03010_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[15\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_98_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07357_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06308_ _00681_ net186 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__nand2_1
XANTENNA__06057__A3 _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07288_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09027_ net251 _04285_ _04287_ net405 net884 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__a32o_1
XFILLER_0_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06239_ net101 _01825_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold250 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[22\]
+ vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[5\]
+ vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[12\] vssd1 vssd1
+ vccd1 vccd1 net942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[11\]
+ vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\] vssd1 vssd1
+ vccd1 vccd1 net964 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout81_A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10870__546 vssd1 vssd1 vccd1 vccd1 _10870__546/HI net546 sky130_fd_sc_hd__conb_1
XANTENNA__05925__A _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10458__RESET_B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09929_ _00701_ _01786_ net155 _04904_ vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__o31a_1
XFILLER_0_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05931__Y _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06756__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06475__B _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10704_ clknet_leaf_68_wb_clk_i _00535_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07493__A2 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ clknet_leaf_44_wb_clk_i _00499_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10566_ clknet_leaf_26_wb_clk_i _00434_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10497_ clknet_leaf_16_wb_clk_i _00365_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10290__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06205__B1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__Y _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput7 wb_rst_i vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07181__A1 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05610_ net445 net444 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__or2_1
X_06590_ net124 _01654_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05541_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] vssd1 vssd1 vccd1
+ vccd1 _01254_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06385__B _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08260_ _03737_ _03738_ net486 vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__o21ba_1
X_05472_ _01059_ _01088_ _01068_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07211_ _02138_ net81 _02750_ _02861_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10338__D team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08191_ _03658_ _03666_ _03669_ _03630_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07142_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[2\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\]
+ net449 vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06444__B1 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07073_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[0\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[8\]
+ net449 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05729__B _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06024_ net197 net205 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__nand2_2
XFILLER_0_61_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10783__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07975_ _03346_ _03432_ _03528_ _03529_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__or4_1
X_09714_ _04733_ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__nor2_1
X_06926_ net433 net150 _02581_ _02501_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09645_ _04705_ _04706_ _04707_ _04708_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__or4_2
X_06857_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout171_X net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05808_ _01494_ _01499_ _01500_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__nor3_1
X_09576_ _04637_ _04661_ net480 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06788_ _01626_ _02412_ _02459_ _01636_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_26_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05480__A _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] _03980_ _03985_
+ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05739_ net1127 _00791_ _01441_ _00766_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[3\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08458_ _03877_ _03930_ net491 net463 _03858_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_136_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07409_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] _02998_
+ net233 vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08389_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] vssd1 vssd1 vccd1
+ vccd1 _03864_ sky130_fd_sc_hd__a21oi_1
X_10420_ clknet_leaf_53_wb_clk_i _00311_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07227__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05238__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10351_ clknet_leaf_40_wb_clk_i _00291_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10282_ clknet_leaf_84_wb_clk_i _00274_ net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_104_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout84_X net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08031__A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09561__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07466__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06674__B1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07218__A2 _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10618_ clknet_leaf_49_wb_clk_i _00482_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07110__A _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06426__B1 _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10549_ clknet_leaf_19_wb_clk_i _00417_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10957__598 vssd1 vssd1 vccd1 vccd1 _10957__598/HI net598 sky130_fd_sc_hd__conb_1
XANTENNA__10244__Q team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06729__A1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__B1 _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ _01067_ net219 net200 _01078_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__o22a_1
XANTENNA__05284__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04972_ net489 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
X_06711_ _02260_ _02262_ _02379_ _02383_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07691_ _01726_ _02365_ _03150_ _01712_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09430_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\]
+ _04577_ _04580_ _04568_ _04579_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06642_ _02108_ _02209_ _02289_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a21o_1
XANTENNA__06396__A _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04909__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09361_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__inv_2
X_06573_ _01687_ _01690_ _02049_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_59_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08312_ _00731_ _01303_ _03677_ _00732_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__o211a_1
X_05524_ _01220_ _01232_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__nand2_1
X_09292_ net228 _04480_ _04482_ net402 net861 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07457__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_12 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ net485 net416 _03721_ net489 vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__a211oi_1
X_05455_ _01156_ _01157_ _01158_ _01159_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_34 team_07_WB.instance_to_wrap.team_07.recFLAG.flagDetect vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout131_A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08174_ _03628_ _03648_ _03634_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05386_ net193 _01000_ _01021_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__nor3_2
XFILLER_0_43_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06562__C _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06417__B1 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07125_ net98 _01616_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07056_ _02688_ _02710_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06007_ net145 net136 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_58_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07958_ _03509_ _03511_ _03512_ _03461_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__a211o_1
XANTENNA__05943__A2 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06909_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] net160 vssd1 vssd1
+ vccd1 vccd1 _02580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07889_ _03443_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__inv_2
X_09628_ _04695_ _04696_ vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_104_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06353__C1 _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09559_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ net800 net236 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09986__RESET_B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06120__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06753__B net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10403_ clknet_leaf_10_wb_clk_i net678 net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09556__S net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ clknet_leaf_51_wb_clk_i net700 net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10876__552 vssd1 vssd1 vccd1 vccd1 _10876__552/HI net552 sky130_fd_sc_hd__conb_1
XFILLER_0_108_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10265_ clknet_leaf_74_wb_clk_i _00257_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10196_ clknet_leaf_84_wb_clk_i _00200_ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05934__A2 _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout390 net392 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05391__Y _01104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06344__C1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07105__A _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06944__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05240_ net302 _00951_ _00952_ vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput10 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput32 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput43 wbs_we_i vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05171_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\]
+ _00883_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07611__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ net436 net867 net244 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08861_ net240 _04191_ _01748_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__o21a_1
XANTENNA__06178__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07812_ _03365_ _03366_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__or2_1
X_08792_ net1026 _04147_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__nand2_1
X_07743_ _03282_ _03287_ _03295_ _03297_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__a22o_1
X_04955_ net434 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XANTENNA__07127__A1 _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout179_A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ _02055_ _02282_ _03227_ _03231_ _01690_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_95_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07015__A _02671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09413_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _02965_ _04557_ _02964_
+ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__a2bb2o_1
X_06625_ _02031_ _02119_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout346_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09344_ net227 _04517_ _04518_ net412 net1095 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06556_ _02229_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05507_ _01219_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
X_09275_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ net1 net337 _04470_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07669__B _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06487_ _02039_ _02042_ _02152_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout134_X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ net4 net3 vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05438_ _00966_ net299 _01136_ _01150_ vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_105_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08157_ net470 net473 vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05369_ _01079_ _01081_ _01078_ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07108_ net159 _01688_ net164 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08088_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[8\]
+ _00814_ net483 vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07039_ _02164_ _02362_ _02184_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05917__B _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09355__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ clknet_leaf_29_wb_clk_i _00108_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06574__C1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05933__A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10952_ net593 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10883_ net559 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_14_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06764__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10317_ clknet_leaf_39_wb_clk_i net743 net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_10248_ clknet_leaf_82_wb_clk_i _00240_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06004__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05546__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10179_ clknet_leaf_8_wb_clk_i _00189_ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07109__A1 _01694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06580__A2 _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__B net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06332__A2 _00754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06410_ _02052_ _02083_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07390_ _02987_ net478 _02986_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[2\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_57_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06341_ _01649_ _02011_ _02015_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_33_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06393__B _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09060_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04310_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__o21a_1
X_06272_ _00684_ net458 net201 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08011_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__xor2_1
X_05223_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00936_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07045__B1 _02699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05154_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[20\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00867_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10972__613 vssd1 vssd1 vccd1 vccd1 _10972__613/HI net613 sky130_fd_sc_hd__conb_1
XANTENNA__07596__A1 _02082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08793__B1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07596__B2 _02744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05085_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00810_ vssd1 vssd1 vccd1
+ vccd1 _00811_ sky130_fd_sc_hd__nand2_1
X_09962_ clknet_leaf_0_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[39\]
+ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08913_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09893_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\] _01775_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout296_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10432__Q team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08844_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\]
+ _04143_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_51_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06849__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06020__A1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08775_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] net711 net245 vssd1
+ vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__mux2_1
X_05987_ net131 net126 _01676_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__and3_2
XFILLER_0_19_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout463_A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ net109 _03280_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__or2_1
X_04938_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] vssd1
+ vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
X_07657_ _03204_ _03214_ _03205_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06608_ _02268_ _02272_ _02273_ _02280_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__o22a_1
X_07588_ _01739_ _03078_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09327_ net228 _04506_ _04507_ net402 net895 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__a32o_1
X_06539_ net119 _02212_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09258_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ _04454_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08209_ net421 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] vssd1 vssd1 vccd1 vccd1
+ _03688_ sky130_fd_sc_hd__and3b_1
X_09189_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05928__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07587__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10102_ clknet_leaf_5_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.displayDetect
+ net317 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.displayPixel
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_112_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10033_ _00053_ _00644_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06759__A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06011__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__D1 _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10935_ net585 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__07511__A1 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10866_ net542 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_38_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10925__670 vssd1 vssd1 vccd1 vccd1 net670 _10925__670/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_30_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10797_ clknet_leaf_77_wb_clk_i _00618_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08775__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07578__A1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06660__C _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05910_ _01583_ net122 _01602_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a21o_2
X_06890_ _02482_ _02560_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05841_ _01524_ _01525_ _01529_ _01522_ _01521_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__a32o_1
XFILLER_0_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08560_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[10\]
+ _03613_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__xor2_1
X_05772_ _01463_ _01470_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07511_ net92 _01609_ _01626_ net100 vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__a31o_1
X_08491_ net140 _03960_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__nand2_2
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07442_ _03019_ _03020_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[21\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07373_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\]
+ _02969_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09112_ net213 _04349_ _04351_ net400 net1112 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__a32o_1
X_06324_ net438 _01396_ net256 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09043_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ _04294_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06255_ net217 _01926_ _01929_ net198 _01930_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__o221a_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05206_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00919_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10822__498 vssd1 vssd1 vccd1 vccd1 _10822__498/HI net498 sky130_fd_sc_hd__conb_1
XFILLER_0_5_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold410 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06186_ _01856_ _01857_ _01863_ _01866_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__o22a_1
XFILLER_0_41_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold421 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[2\] vssd1
+ vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold443 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\] vssd1 vssd1
+ vccd1 vccd1 net1113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__dlygate4sd3_1
X_05137_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00850_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold465 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\] vssd1 vssd1 vccd1
+ vccd1 net1135 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\] vssd1 vssd1
+ vccd1 vccd1 net1146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 team_07_WB.instance_to_wrap.team_07.label_num_bus\[26\] vssd1 vssd1 vccd1
+ vccd1 net1157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\] vssd1 vssd1
+ vccd1 vccd1 net1168 sky130_fd_sc_hd__dlygate4sd3_1
X_05068_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back _00795_
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select vssd1
+ vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__or4b_4
XFILLER_0_110_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09945_ net463 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ net964 _04871_ _04872_ vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__o21a_1
X_08827_ _04171_ _04172_ net195 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07741__A1 _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08758_ net944 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ net239 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07709_ net156 net202 net172 _01744_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__o31a_1
XFILLER_0_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08689_ _00707_ _04105_ _04108_ _04110_ vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__o31a_1
XFILLER_0_135_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ clknet_leaf_62_wb_clk_i _00551_ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05930__B net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10651_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_sck_fl_enable
+ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.sck_fl_enable
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10246__RESET_B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10582_ clknet_leaf_53_wb_clk_i _00446_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_106_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09549__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09564__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__A1 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ clknet_leaf_43_wb_clk_i net899 net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06639__D net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06001__B net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10918_ net663 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_128_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08693__C1 _01759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10849_ net525 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
XFILLER_0_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08445__C1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06952__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07767__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06671__B _02027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06040_ _01668_ _01715_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__or2_2
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06016__X _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout208 net209 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout219 _01502_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_8
X_07991_ net259 _03437_ _03450_ _03505_ _03545_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recGen.circleDetect
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_10_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09730_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06942_ _02500_ _02509_ net201 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__a21oi_1
XANTENNA__05982__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06399__A net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09661_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\] _04720_ vssd1
+ vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__and2_1
XANTENNA__07478__C_N _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06873_ _02466_ _02474_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__or2_1
XANTENNA__06526__A2 _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08612_ _01109_ _01926_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__nand2_1
X_05824_ _01513_ _01516_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__nand2_1
X_09592_ _04665_ _04672_ _04669_ net1039 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08543_ _03608_ _03995_ _03999_ vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__a21oi_1
X_05755_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[24\] vssd1 vssd1 vccd1
+ vccd1 _01454_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout161_A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout259_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05686_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[0\] net440 vssd1 vssd1
+ vccd1 vccd1 _01399_ sky130_fd_sc_hd__or2_1
X_08474_ _03911_ _03930_ _03945_ net415 vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07425_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\] _03008_
+ net478 vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10936__X net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07356_ net477 _02963_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_21_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06307_ net187 _01975_ _01982_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_135_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07287_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09026_ _04286_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06462__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06238_ _01888_ _01910_ _01916_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simonGen.simonDetect\[2\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06169_ _01849_ _01809_ _01817_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__and3b_1
Xhold240 _00467_ vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[33\]
+ vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[0\] vssd1
+ vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07693__A _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07411__B1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 _00099_ vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[3\] vssd1 vssd1
+ vccd1 vccd1 net965 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09928_ net340 _01785_ _01790_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\]
+ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09859_ _04666_ _04731_ _04767_ net269 team_07_WB.instance_to_wrap.audio vssd1 vssd1
+ vccd1 vccd1 _04861_ sky130_fd_sc_hd__o41a_1
XFILLER_0_99_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05941__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10703_ clknet_leaf_68_wb_clk_i _00534_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05899__B1_N _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09559__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10634_ clknet_leaf_44_wb_clk_i net840 net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10565_ clknet_leaf_26_wb_clk_i _00433_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06491__B net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10496_ clknet_leaf_15_wb_clk_i _00364_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output55_A net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08902__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05540_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__nor2_1
XANTENNA__07469__B1 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06385__C net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05471_ _01034_ _01080_ _01183_ _01145_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__o31a_1
XFILLER_0_117_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07210_ _02856_ _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__or2_1
X_08190_ _03631_ _03668_ _00717_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__mux2_1
XANTENNA__06692__A1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06682__A _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07141_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] net301 net300 team_07_WB.instance_to_wrap.team_07.label_num_bus\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07072_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\] _00831_ _00942_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[25\]
+ _02725_ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06023_ net1133 _01633_ _01641_ _01713_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[2\]
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_26_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07974_ _03340_ _03425_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09713_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\] net250 _04754_
+ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__and3_1
X_06925_ _02593_ _02595_ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__nor2_1
X_09644_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__or4b_1
XANTENNA__10591__RESET_B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06856_ _02475_ _02492_ _02493_ _02526_ _01689_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a2111o_1
XANTENNA__06857__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05807_ _01499_ _01500_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__nor2_1
X_09575_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] _04661_
+ _04662_ vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__a21bo_1
X_06787_ _00674_ _02332_ _02170_ net431 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a211oi_1
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _03980_ _03985_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05480__B _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05738_ _00652_ _00773_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08457_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[0\] _03744_ _03804_
+ _03929_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__or4_1
XANTENNA__06132__B1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05669_ _01381_ vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07408_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] _02998_
+ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ net794 net130 _03832_ _03863_ vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07339_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ _02411_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09621__A1 _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07227__A3 _02276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05238__A2 team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10350_ clknet_leaf_40_wb_clk_i _00290_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09009_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10281_ clknet_leaf_0_wb_clk_i _00273_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05936__A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08031__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05942__Y _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__A2 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06123__B1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06674__A1 _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10617_ clknet_leaf_49_wb_clk_i _00481_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07110__B _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548_ clknet_leaf_19_wb_clk_i _00416_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06007__A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479_ clknet_leaf_22_wb_clk_i _00347_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04971_ net418 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
X_06710_ _02154_ _02260_ _02382_ _02381_ _02380_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a32o_1
XFILLER_0_95_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07690_ _01631_ _02009_ _02348_ net94 net100 vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__o221a_1
XANTENNA__05581__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06641_ _00635_ _02212_ _02305_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06396__B _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ _04525_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__and3_1
X_06572_ net204 _02066_ _02171_ _02164_ _02158_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10600__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08103__A1 _03604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08311_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\] _01308_ _01384_
+ _03788_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[3\] vssd1 vssd1
+ vccd1 vccd1 _03789_ sky130_fd_sc_hd__a311o_1
X_05523_ _01220_ _01232_ _01235_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__o22a_1
X_09291_ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__inv_2
XANTENNA__06114__B1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_13 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _03672_ _03720_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__nor2_1
X_05454_ net299 _01029_ _01092_ _01154_ _01155_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_24 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_59_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08173_ _03628_ _03648_ _03634_ vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__a21o_1
X_05385_ _01096_ _01097_ _01094_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_132_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout124_A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06417__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ _02729_ _02763_ _02777_ _01646_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10435__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07055_ _02681_ _02677_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06006_ net148 net132 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__nor2_8
XFILLER_0_11_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07917__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__B2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10772__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ _03288_ _03391_ _03351_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06908_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] _01557_ vssd1 vssd1
+ vccd1 vccd1 _02579_ sky130_fd_sc_hd__or2_1
X_07888_ _01078_ net161 vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__nand2_1
X_09627_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[16\] _04694_ vssd1
+ vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__and2_1
X_06839_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] _02498_ _02509_
+ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__o21ai_2
XANTENNA__06353__B1 _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09558_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ net796 net236 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08509_ _03969_ _03970_ _03972_ _03973_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09489_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[17\]
+ net270 _04619_ net290 net220 vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10402_ clknet_leaf_10_wb_clk_i net692 net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08948__A3 _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10333_ clknet_leaf_51_wb_clk_i net707 net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_10264_ clknet_leaf_74_wb_clk_i _00256_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10195_ clknet_leaf_90_wb_clk_i _00199_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05953__X _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10080__Q net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_2
XANTENNA__05934__A3 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06895__A1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08097__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput11 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput22 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput33 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05170_ _00849_ _00877_ _00882_ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07775__B net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08860_ _00797_ _00959_ _00960_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__nor3_1
X_07811_ _01095_ net147 vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_88_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08791_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\] _04147_ vssd1
+ vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__or2_1
X_07742_ _03281_ _03283_ _03296_ _03276_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_79_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04954_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1 vssd1 vccd1
+ vccd1 _00694_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07127__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07673_ net156 _03229_ _03230_ _03228_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__a211o_1
XANTENNA__06335__B1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09412_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _02965_ _04556_ _02963_
+ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__o22a_2
X_06624_ _02285_ _02294_ _02296_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09343_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ _04514_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__or2_1
XANTENNA__08088__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06555_ net157 _01644_ net202 _01663_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout339_A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05506_ _01207_ _01217_ _01218_ net422 net424 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__o32a_1
X_09274_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ net1 _04263_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06486_ _02092_ _02155_ _02153_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08225_ net5 _03703_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__and2b_1
X_05437_ _01130_ _01148_ _01149_ _01136_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__or4b_1
XANTENNA__10944__X net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout127_X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08156_ net470 net473 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nor2_2
X_05368_ _01080_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07063__A1 _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ net82 _02759_ _02760_ net98 _01635_ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__o221a_4
XFILLER_0_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08087_ _03596_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[8\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__mux2_1
X_05299_ _01009_ _01011_ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__nand2_1
X_07038_ _02692_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08989_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__and3_1
XANTENNA__06574__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05933__B _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10951_ net592 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_123_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06877__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10882_ net558 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_97_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07212__Y _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05852__A2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07054__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10694__RESET_B net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05396__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10316_ clknet_leaf_39_wb_clk_i net746 net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10247_ clknet_leaf_82_wb_clk_i _00239_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06004__B net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07498__A_N _00943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ clknet_leaf_9_wb_clk_i _00188_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10930__580 vssd1 vssd1 vccd1 vccd1 _10930__580/HI net580 sky130_fd_sc_hd__conb_1
XANTENNA__06580__A3 _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08857__A2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06332__A3 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06340_ _01723_ _02012_ _02013_ net418 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06271_ net183 _01929_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05222_ _00933_ _00934_ _00932_ vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__a21oi_1
X_08010_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06690__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05153_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__and2b_1
XANTENNA__07045__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05084_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\] _00808_
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\] vssd1
+ vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__and4bb_1
X_09961_ clknet_leaf_85_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[38\]
+ net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06715__A_N _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08912_ net264 _04221_ vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09892_ net1093 net154 net152 _04882_ vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__a22o_1
X_08843_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\] _04143_
+ net908 vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_51_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06020__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] net687 net245 vssd1
+ vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05986_ net133 net129 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__nand2_8
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07725_ _03273_ _03274_ _03275_ _03278_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_0_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04937_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\] vssd1
+ vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
XANTENNA__08848__A2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06859__A1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ net144 _01689_ _01730_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__or3_1
XANTENNA__06859__B2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06865__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10827__503 vssd1 vssd1 vccd1 vccd1 _10827__503/HI net503 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_74_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_06607_ _02266_ _02274_ _02279_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__and3b_1
XFILLER_0_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07587_ net187 net106 net142 _01671_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout244_X net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05531__B2 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09326_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ _04502_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__nand3_1
XFILLER_0_75_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06538_ net288 _01620_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__or2_2
XFILLER_0_36_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09257_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ _04454_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06469_ _02068_ _02101_ _02105_ _02107_ _02130_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07696__A _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08208_ _01261_ _03686_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__nand2_1
X_09188_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ _04404_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08139_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[23\] _03623_
+ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_116_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05928__B net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07587__A2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05647__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ clknet_leaf_31_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.buttonDetect
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.buttonPixel sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05944__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10032_ _00052_ _00643_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__06011__A2 _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10934_ net584 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07511__A2 _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10865_ net541 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ clknet_leaf_78_wb_clk_i _00617_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10995__636 vssd1 vssd1 vccd1 vccd1 _10995__636/HI net636 sky130_fd_sc_hd__conb_1
XFILLER_0_22_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06015__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05557__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06786__A0 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06002__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05840_ _00714_ _01530_ _01533_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_55_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05771_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\] _01469_
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\]
+ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__and4bb_1
X_07510_ _03066_ _03067_ _03068_ _03065_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__o31a_1
X_08490_ _03633_ _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07441_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] _03018_
+ _02984_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10341__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07372_ _02974_ _02975_ _02976_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[2\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07634__B1_N _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09111_ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06323_ _01972_ _01991_ _01994_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09042_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ _04291_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__a31o_1
X_06254_ net458 net217 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05205_ _00916_ _00917_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_96_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold400 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.next_back vssd1
+ vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06185_ _01856_ _01865_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__nand2b_1
Xhold411 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[0\] vssd1 vssd1 vccd1
+ vccd1 net1081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\] vssd1 vssd1
+ vccd1 vccd1 net1092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\] vssd1 vssd1
+ vccd1 vccd1 net1103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05136_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__nor2_1
Xhold444 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] vssd1 vssd1
+ vccd1 vccd1 net1114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06777__B1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold466 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 net52 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold488 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05067_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back _00795_
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select vssd1
+ vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__nor4b_4
X_09944_ net463 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
Xhold499 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[0\] vssd1
+ vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08019__A_N net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08778__C net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ net153 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__or3b_1
XANTENNA_input9_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08826_ net1115 _04141_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__nand2_1
XANTENNA__07741__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08757_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[31\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ net235 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__mux2_1
X_05969_ net255 _01658_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07708_ _01675_ _03261_ _03262_ _03263_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08688_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ net457 _04073_ _04107_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__a41o_1
XANTENNA__06595__A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _01655_ _01728_ _01874_ _03196_ net260 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a2111o_1
XANTENNA__05930__C _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10650_ clknet_leaf_40_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_sck_rs_enable
+ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.sck_rs_enable
+ sky130_fd_sc_hd__dfrtp_1
X_09309_ _04494_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10581_ clknet_leaf_62_wb_clk_i _00012_ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_118_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10286__RESET_B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06106__Y _01789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05945__Y _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05991__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ clknet_leaf_43_wb_clk_i _00094_ net387 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09433__X _04582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06001__C _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10917_ net662 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10848_ net524 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_67_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10779_ clknet_leaf_65_wb_clk_i _00600_ net356 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06671__C _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07956__C1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout209 _04583_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_4
X_07990_ _03532_ _03537_ _03538_ _03544_ _03531_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06941_ net433 _02500_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] vssd1
+ vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
XANTENNA__05982__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06399__B _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09660_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\]
+ _04717_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06872_ net434 _02528_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__nor2_1
X_08611_ _04041_ _04040_ _04037_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_59_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05823_ _01513_ _01516_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__and2_1
X_09591_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ _04671_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ _03996_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05754_ _01448_ _01451_ _01452_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__or3_1
XANTENNA__04928__A team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08473_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\] _03944_
+ _03713_ net465 vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__o211a_1
X_05685_ net441 net440 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_46_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07424_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\] _03008_
+ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07239__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07355_ _02963_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout321_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06306_ _01974_ _01976_ _01981_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_135_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07286_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__nor2_1
X_09025_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ _04280_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06462__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06237_ _01838_ _01869_ _01875_ _01915_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__and4b_1
XFILLER_0_115_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold230 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__dlygate4sd3_1
X_06168_ net289 _01679_ _01689_ _01848_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a31o_1
Xhold241 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[4\]
+ vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[32\]
+ vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[43\]
+ vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__dlygate4sd3_1
X_05119_ net302 _00830_ vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__nor2_1
Xhold274 team_07_WB.instance_to_wrap.team_07.label_num_bus\[32\] vssd1 vssd1 vccd1
+ vccd1 net944 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07693__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold285 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[13\]
+ vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__dlygate4sd3_1
X_06099_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[17\]
+ _01781_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__or3_1
Xhold296 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\] vssd1 vssd1
+ vccd1 vccd1 net966 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09927_ _01785_ net151 _04903_ net838 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09858_ net1120 _04824_ _04860_ _04805_ vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08809_ net969 _04160_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09789_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\] _04808_ _04812_
+ vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__a21o_1
XANTENNA__05941__B net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10702_ clknet_leaf_68_wb_clk_i _00533_ net347 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06150__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10633_ clknet_leaf_48_wb_clk_i _00497_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10564_ clknet_leaf_26_wb_clk_i _00432_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06491__C net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10495_ clknet_leaf_16_wb_clk_i _00363_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07108__B _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10414__SET_B net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09458__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07469__A1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05470_ _01061_ _01096_ _01064_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06141__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06692__A2 _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07140_ _02791_ _02792_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_41_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07071_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[33\] net302 net398 _02724_
+ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06022_ net144 _01667_ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__nand2_2
XANTENNA__07794__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06601__C1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07973_ _03525_ _03527_ _03526_ _03367_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__or4b_1
X_09712_ _04754_ _04755_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\]
+ _04730_ vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__a2bb2o_1
X_06924_ net174 _02511_ _02594_ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__o21ai_1
X_09643_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__nand4b_1
X_06855_ _02525_ _02503_ _02497_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout271_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout369_A net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05806_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\] _01496_
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] vssd1 vssd1
+ vccd1 vccd1 _01500_ sky130_fd_sc_hd__and3b_1
X_09574_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] _01418_
+ _04661_ net480 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__o31a_1
XANTENNA__06380__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06786_ net431 _02413_ _00673_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__mux2_1
X_08525_ net987 _03978_ _03986_ vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07034__A _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05737_ _01437_ _01440_ _01439_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[1\]
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_65_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout157_X net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08456_ _03709_ _03928_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_137_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06132__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05668_ _00678_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] vssd1 vssd1 vccd1
+ vccd1 _01381_ sky130_fd_sc_hd__nor3_2
XFILLER_0_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07407_ _02998_ net233 _02997_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[8\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_136_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08387_ _03753_ _03862_ _03653_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07880__A1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06592__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05599_ _01305_ _01306_ _01311_ vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07338_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[2\] team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07269_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ _02904_ _02907_ _01315_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[17\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_130_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09008_ net251 _04272_ _04273_ net403 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__a32o_1
XFILLER_0_103_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10280_ clknet_leaf_87_wb_clk_i _00272_ net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05936__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05946__A1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07148__B1 _02781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05952__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10648__RESET_B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06123__A1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08327__X _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06674__A2 _01582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10616_ clknet_leaf_49_wb_clk_i _00480_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10547_ clknet_leaf_19_wb_clk_i _00415_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07623__A1 _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06007__B net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10478_ clknet_leaf_22_wb_clk_i _00346_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09318__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__A2 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_04970_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row vssd1 vssd1 vccd1
+ vccd1 _00709_ sky130_fd_sc_hd__inv_2
X_06640_ _02312_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06571_ _02129_ _02242_ _02243_ _02244_ _02241_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_87_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08310_ _01306_ _03682_ _03786_ _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__o211a_1
X_05522_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ _01232_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__nor2_1
X_09290_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ _04475_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06114__A1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06693__A _02209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08241_ team_07_WB.instance_to_wrap.team_07.circlePixel net485 vssd1 vssd1 vccd1
+ vccd1 _03720_ sky130_fd_sc_hd__nand2b_1
XANTENNA__06665__A2 _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_14 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07862__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05453_ _01057_ _01075_ _01111_ _01160_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_60_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_25 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07862__B2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860__536 vssd1 vssd1 vccd1 vccd1 _10860__536/HI net536 sky130_fd_sc_hd__conb_1
XFILLER_0_16_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08172_ _03628_ _03648_ _03651_ _03649_ net466 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__a32o_1
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05384_ net194 _01005_ _01021_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_132_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07123_ _02764_ _02767_ _02776_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07614__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06417__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07054_ net276 net274 _01638_ _02335_ _02708_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__o311a_1
XANTENNA__08413__A _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06005_ net158 net147 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__or2_4
XFILLER_0_101_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_28_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_58_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10451__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ _01057_ _01741_ _03371_ _03510_ net256 vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__o221a_1
X_06907_ net433 net182 _02505_ _02577_ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a211o_1
XANTENNA__08878__B1 _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07887_ _01078_ net161 vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06587__B _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09626_ net1072 _04694_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__nor2_1
X_06838_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__nand2_2
XANTENNA__06353__A1 _00709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09557_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ net721 net236 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__mux2_1
X_06769_ _02417_ _02440_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__nor2_1
X_08508_ _03969_ _03970_ _03972_ _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07699__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09488_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _04616_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_121_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08439_ net462 _03912_ _03681_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05012__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10401_ clknet_leaf_9_wb_clk_i net686 net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_116_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07605__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ clknet_leaf_52_wb_clk_i net701 net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10263_ clknet_leaf_74_wb_clk_i _00255_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10194_ clknet_leaf_84_wb_clk_i _00198_ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout370 net375 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_4
Xfanout381 net388 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_2
Xfanout392 net75 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10411__RESET_B net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05855__B1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput12 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput34 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07057__C1 _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07810_ _01094_ net145 vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_88_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05863__Y _01557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08790_ _04147_ _04148_ net196 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_88_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05592__A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07741_ _01064_ net117 _03291_ _00750_ _03290_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__o221a_1
XANTENNA__06040__X _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04953_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07672_ _01680_ _02055_ _02081_ _01646_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__a22o_1
XANTENNA__06335__A1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07532__B1 _03075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09411_ net857 _04566_ _04565_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__mux2_1
X_06623_ _02280_ _02292_ _02269_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a21o_1
XANTENNA__10598__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09342_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ _04514_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__nand2_1
X_06554_ _02139_ net85 _02214_ _02149_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05505_ _01199_ _01216_ _01210_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09273_ net3 net1185 _04469_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06485_ _01636_ _02157_ _02158_ _02109_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ net6 net1 vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05436_ net435 _01072_ _01131_ net299 _01146_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10899__565 vssd1 vssd1 vccd1 vccd1 _10899__565/HI net565 sky130_fd_sc_hd__conb_1
X_08155_ net470 net472 vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout401_A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05367_ net191 _01025_ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__nor2_1
X_07106_ _01630_ _01636_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08086_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[7\]
+ _00814_ net483 vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__o21a_1
XANTENNA__07063__A2 _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05298_ net192 _01004_ _01010_ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07037_ _02677_ _02681_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_77_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06023__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08988_ net2 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ _04257_ vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07939_ _01078_ net200 net189 _01084_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_3_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10950_ net591 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_123_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06326__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07523__B1 _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09609_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\] _04682_ vssd1
+ vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__or2_1
X_10881_ net557 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_79_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10947__588 vssd1 vssd1 vccd1 vccd1 _10947__588/HI net588 sky130_fd_sc_hd__conb_1
XANTENNA__07222__A _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08037__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05948__Y _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07054__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10315_ clknet_leaf_39_wb_clk_i net775 net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10246_ clknet_leaf_76_wb_clk_i _00238_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_10177_ clknet_leaf_9_wb_clk_i _00187_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07109__A3 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07132__A _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06270_ net138 _01926_ _01928_ net159 _01946_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05221_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00934_ sky130_fd_sc_hd__or2_1
XANTENNA__06690__B _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05152_ _00861_ _00864_ vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05083_ _00705_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\] vssd1
+ vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__or3_1
X_09960_ clknet_leaf_90_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[29\]
+ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08911_ net438 _01400_ _01403_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__a31o_1
X_09891_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\] _01775_ vssd1
+ vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08568__A_N net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08842_ net976 _04143_ _04181_ vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_51_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07307__A _02930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08773_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] net690 net245 vssd1
+ vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__mux2_1
XANTENNA__06020__A3 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05985_ net135 net125 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__nor2_8
XFILLER_0_109_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout184_A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07724_ _03273_ _03278_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04936_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\] vssd1 vssd1
+ vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07505__B1 _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07655_ _02734_ _03181_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout351_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10866__542 vssd1 vssd1 vccd1 vccd1 _10866__542/HI net542 sky130_fd_sc_hd__conb_1
XANTENNA_fanout449_A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ net134 net127 _01936_ _02275_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__or4_1
X_07586_ net260 net184 _02151_ _01663_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__o31a_1
XFILLER_0_94_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09325_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ _04499_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__a31o_1
XANTENNA__07042__A _02086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06537_ _02208_ _02210_ _02207_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09256_ net230 _04456_ _04457_ net406 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06468_ _02119_ _02126_ _02133_ _01625_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06881__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08207_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] _03682_
+ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__nor2_1
XANTENNA__06492__B1 _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05419_ _01034_ _01036_ _01039_ _01099_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__or4_1
Xclkbuf_leaf_43_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09187_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ _04404_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__or2_1
XANTENNA__07696__B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06399_ net175 _01732_ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__nand2_4
XFILLER_0_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08138_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[23\]
+ _03624_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07587__A3 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[0\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10100_ clknet_leaf_31_wb_clk_i team_07_WB.instance_to_wrap.team_07.memGen.stageDetect
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.stagePixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08601__A team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _00051_ _00047_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05944__B net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10933_ net583 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07511__A3 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ net540 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_67_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10795_ clknet_leaf_77_wb_clk_i _00616_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05959__X _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07887__A _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06483__B1 _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06015__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10229_ clknet_leaf_0_wb_clk_i _00233_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08230__B team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06031__A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05770_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[9\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] vssd1 vssd1 vccd1
+ vccd1 _01469_ sky130_fd_sc_hd__nand3_1
XFILLER_0_89_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07440_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\] _03018_
+ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06710__A1 _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07371_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\] _02969_
+ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09110_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ _04347_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__and2_1
X_06322_ _01972_ _01983_ _01994_ _01997_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09041_ net252 _04296_ _04297_ net407 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__a32o_1
XFILLER_0_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06253_ net217 _01926_ _01929_ net198 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05204_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00917_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold401 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\] vssd1 vssd1
+ vccd1 vccd1 net1071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06184_ net175 net120 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__xnor2_1
Xhold412 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold423 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\] vssd1 vssd1
+ vccd1 vccd1 net1093 sky130_fd_sc_hd__dlygate4sd3_1
X_05135_ _00845_ _00847_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold434 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] vssd1 vssd1
+ vccd1 vccd1 net1115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold456 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__dlygate4sd3_1
X_05066_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ _00793_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__or2_2
Xhold489 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\] vssd1
+ vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ net463 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_wb_clk_i_X clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ net983 net153 _04871_ vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__a21o_1
XANTENNA__06529__A1 _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[16\] _04141_
+ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout187_X net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06544__A4 _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08756_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[30\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[30\]
+ net234 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__mux2_1
X_05968_ net255 net218 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__nand2_1
X_04919_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
X_07707_ _02040_ _02877_ _01744_ _01795_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__a211o_1
X_08687_ _04046_ _04109_ vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__nor2_1
X_05899_ _01591_ _01592_ _01574_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_36_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07638_ _01644_ _01675_ _01742_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_68_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07569_ _01611_ _02332_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09308_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ _04491_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10580_ clknet_leaf_61_wb_clk_i _00011_ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09239_ net231 _04443_ _04445_ net408 net783 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06116__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05020__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06768__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05955__A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10149__SET_B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05991__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ clknet_leaf_42_wb_clk_i net957 net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05961__Y _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10962__603 vssd1 vssd1 vccd1 vccd1 _10962__603/HI net603 sky130_fd_sc_hd__conb_1
X_10916_ net661 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_0_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08693__A1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09890__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ net523 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_39_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08445__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10778_ clknet_leaf_65_wb_clk_i _00599_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06456__B1 _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06026__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06940_ _02522_ _02596_ _02605_ _02610_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06032__Y _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05982__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06871_ _02533_ _02541_ net136 _02526_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08610_ _00689_ _01201_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05822_ _01492_ _01493_ _01501_ _01515_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__o31a_2
X_09590_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\] vssd1 vssd1 vccd1 vccd1
+ _04671_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06931__B2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08541_ _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__inv_2
X_05753_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[14\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\] vssd1 vssd1 vccd1
+ vccd1 _01452_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08472_ _03770_ _03942_ _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05684_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[0\] team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07423_ _03008_ net478 _03007_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[14\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout147_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07354_ _02961_ _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_98_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07239__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06305_ _01978_ _01979_ _01980_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__and3b_1
XFILLER_0_115_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07285_ net1184 _02914_ _02917_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[11\]
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_135_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ _04283_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06236_ net101 _01671_ _01874_ _01914_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold220 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06167_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] net127
+ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__xnor2_1
Xhold231 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout102_X net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[14\]
+ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__dlygate4sd3_1
X_05118_ net450 team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\] _00685_ vssd1
+ vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__and3b_1
Xhold264 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[12\]
+ vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__dlygate4sd3_1
X_06098_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[15\] _01780_
+ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__or2_1
Xhold275 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[9\]
+ vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[5\]
+ vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09926_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\] _01784_
+ net155 vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__or3_1
X_05049_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00780_ vssd1 vssd1
+ vccd1 vccd1 _00781_ sky130_fd_sc_hd__nand2_1
X_10915__660 vssd1 vssd1 vccd1 vccd1 net660 _10915__660/LO sky130_fd_sc_hd__conb_1
X_09857_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[15\] _04858_ vssd1
+ vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08808_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\] _04154_ vssd1 vssd1
+ vccd1 vccd1 _04160_ sky130_fd_sc_hd__or4_2
X_09788_ _01768_ _04810_ _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08739_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ net234 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10701_ clknet_leaf_68_wb_clk_i _00532_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06150__A2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10632_ clknet_leaf_49_wb_clk_i _00496_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10563_ clknet_leaf_24_wb_clk_i _00431_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05021__Y _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07650__A2 _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10494_ clknet_leaf_15_wb_clk_i _00362_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06429__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07070_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[1\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[9\]
+ net449 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05298__C _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06021_ net137 _01708_ _01712_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__or3_1
XANTENNA__07794__B _01069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05404__A1 _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07972_ _01113_ net178 net256 vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__o21ai_1
X_09711_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] _04752_ _04731_
+ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__o21ai_1
X_06923_ net190 _02508_ _02577_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07157__A1 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09642_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__or4_1
XFILLER_0_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06854_ _02499_ _02504_ _02524_ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_93_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05805_ _01495_ _01496_ _01498_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__a21oi_2
X_09573_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ _04629_ _04657_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__or3_2
X_06785_ _02410_ _02414_ net94 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06380__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08524_ _03985_ _03976_ _03984_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__or3b_1
X_05736_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ _00652_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08455_ net486 net488 net489 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__or4b_1
X_05667_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] vssd1 vssd1 vccd1
+ vccd1 _01380_ sky130_fd_sc_hd__nor3b_1
XANTENNA_fanout431_A team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06132__A2 _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07406_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\]
+ _02994_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_82_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08386_ net465 _03859_ _03861_ _03749_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__o22a_1
X_05598_ _01303_ _01304_ _01302_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07337_ _02947_ _02949_ _02936_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[1\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07268_ _01315_ _02907_ _02908_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[16\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06219_ net96 _01878_ _01885_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09007_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__nand3_1
XFILLER_0_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07199_ _01739_ _02036_ _02836_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05946__A2 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\] _01779_
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[14\] vssd1 vssd1 vccd1
+ vccd1 _04893_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_109_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05952__B _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08755__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06674__A3 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10615_ clknet_leaf_52_wb_clk_i _00479_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05399__B _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10546_ clknet_leaf_19_wb_clk_i _00414_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07623__A2 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10477_ clknet_leaf_22_wb_clk_i _00345_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06304__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06570_ _02050_ _02114_ _02134_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05521_ _01219_ _01232_ _01233_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06114__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08240_ team_07_WB.instance_to_wrap.team_07.circlePixel net485 vssd1 vssd1 vccd1
+ vccd1 _03719_ sky130_fd_sc_hd__and2b_1
X_05452_ _01163_ _01164_ vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_15 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_26 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10358__RESET_B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08171_ net53 _03628_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__or2_1
X_05383_ _01001_ net192 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07122_ _02768_ _02773_ _02775_ _02277_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06417__A3 _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10901__567 vssd1 vssd1 vccd1 vccd1 _10901__567/HI net567 sky130_fd_sc_hd__conb_1
XFILLER_0_43_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07053_ net86 net253 _01639_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a21o_1
XANTENNA__06283__D1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06004_ net159 net148 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_68_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07955_ net162 _03375_ _03458_ _03462_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout381_A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08327__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ net432 net182 _02517_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_98_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07886_ _01078_ net161 vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__nor2_1
X_09625_ _04664_ _04693_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__nor2_1
X_06837_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07550__A1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout267_X net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06353__A2 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09556_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ net823 net243 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__mux2_1
X_06768_ net431 net276 _02413_ _02439_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08507_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__and4bb_1
X_05719_ net482 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ _00822_ _01429_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_121_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06699_ net258 _02014_ _02048_ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a21o_1
X_09487_ net936 net206 _04618_ vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08438_ _00730_ _01284_ _03689_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__o21a_1
XANTENNA__10099__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08369_ net459 _03842_ _03843_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_34_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ clknet_leaf_10_wb_clk_i net709 net325 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07605__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05616__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10331_ clknet_leaf_52_wb_clk_i net703 net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05439__S _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10262_ clknet_leaf_74_wb_clk_i _00254_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06124__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ clknet_leaf_90_wb_clk_i _00197_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout82_X net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05963__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06411__X _02085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout360 net361 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_4
Xfanout371 net374 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout382 net384 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_4
Xfanout393 _03562_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08869__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06130__Y _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06344__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10883__559 vssd1 vssd1 vccd1 vccd1 _10883__559/HI net559 sky130_fd_sc_hd__conb_1
XFILLER_0_51_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput13 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput24 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput35 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10529_ clknet_leaf_25_wb_clk_i _00397_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06034__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10818__494 vssd1 vssd1 vccd1 vccd1 _10818__494/HI net494 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_88_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04952_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
X_07740_ net268 _03285_ _03294_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__or3_1
XANTENNA__05592__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ net107 _01719_ net165 _01678_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__a22o_1
XANTENNA__06335__A2 _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09410_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _04556_ vssd1 vssd1 vccd1
+ vccd1 _04566_ sky130_fd_sc_hd__nor2_1
X_06622_ _01714_ _01742_ _02294_ _02293_ _02267_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_94_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09341_ net227 _04515_ _04516_ net412 net913 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__a32o_1
X_06553_ _02085_ _02131_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05504_ _01203_ _01211_ _01212_ _01214_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__a31o_1
X_09272_ _04420_ _04422_ _04466_ _04468_ _04421_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__a2111o_1
X_06484_ _02057_ _02155_ _02153_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08223_ _03700_ _03701_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__o21ai_2
X_05435_ _01141_ _01142_ _01143_ _01147_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__or4b_1
XFILLER_0_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07048__B1 _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ net470 net472 vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__and2_1
X_05366_ net194 _01074_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07105_ _01636_ _02197_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__nor2_1
X_08085_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[7\]
+ net232 _03595_ net898 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07063__A3 _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05297_ net431 _00998_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__nand2_2
XFILLER_0_114_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07036_ _02111_ _02687_ _02690_ _02685_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_77_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10462__Q team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08987_ _04250_ _04251_ _04254_ _04256_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__or4_1
X_07938_ _01692_ _03492_ _03490_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09512__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07869_ net282 net397 _01063_ _03350_ _03423_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_123_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07523__A1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09608_ _00697_ _04680_ _04682_ _04665_ vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__a22oi_1
X_10880_ net556 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_94_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09539_ _04650_ net925 net223 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07222__B _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05023__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05958__A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10314_ clknet_leaf_46_wb_clk_i net793 net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_104_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05964__Y _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ clknet_leaf_75_wb_clk_i _00237_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07892__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07237__X _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ clknet_leaf_9_wb_clk_i _00186_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 _01531_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload5_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10632__RESET_B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08228__B _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07132__B _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08475__C1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07700__X _03256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06971__B net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05220_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00933_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06690__C net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05151_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00864_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07045__A3 _02697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06253__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05082_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[1\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[0\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__and3_1
XANTENNA__06253__B2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08910_ net264 _04220_ vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09890_ net841 net153 net151 _04881_ vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08841_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\] _01457_
+ _04143_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08772_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\] net834 net245 vssd1
+ vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__mux2_1
X_05984_ net160 net150 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__or2_4
XFILLER_0_58_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07723_ _01597_ _01604_ _01105_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__a21oi_1
X_04935_ net431 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07505__A1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout177_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07654_ _01730_ _02765_ _03160_ _03211_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__o31ai_1
XANTENNA__04947__A team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06605_ net107 _01935_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__nand2_2
X_07585_ _02107_ _02164_ net87 vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_137_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09324_ net228 _04504_ _04505_ net401 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05114__Y _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06536_ _02178_ _02209_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10907__573 vssd1 vssd1 vccd1 vccd1 _10907__573/HI net573 sky130_fd_sc_hd__conb_1
XFILLER_0_35_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09255_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ _04454_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06467_ _02060_ _02092_ _02090_ _02068_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_90_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05778__A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ _03683_ _03684_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_79_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05418_ _01017_ _01033_ _01041_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__or3_1
X_09186_ net211 _04403_ _04405_ net402 net1056 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__a32o_1
X_06398_ _02071_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__inv_2
XANTENNA__08769__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08137_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ _03623_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__nor2_1
X_05349_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] net436 vssd1
+ vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_116_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08068_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ _03024_ net298 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ _03587_ vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07019_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\]
+ net449 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_12_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10030_ _00050_ _00046_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06402__A _02060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__A1 _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05018__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10932_ net582 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_129_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06294__A1_N net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10863_ net539 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_67_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10794_ clknet_leaf_77_wb_clk_i _00615_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07887__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10438__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07680__B1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07983__B2 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05994__B1 _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10228_ clknet_leaf_85_wb_clk_i _00232_ net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06312__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__A0 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10159_ clknet_leaf_3_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[6\]
+ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold2 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06031__B _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08239__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06710__A2 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07370_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\] _02969_
+ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06321_ _01981_ _01996_ _01995_ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07797__B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09040_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ _04294_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06252_ _01926_ _01927_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__nand2_2
XANTENNA__07671__B1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05203_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00916_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06183_ net175 net120 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_96_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold402 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[16\] vssd1 vssd1
+ vccd1 vccd1 net1072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold413 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[11\] vssd1 vssd1
+ vccd1 vccd1 net1083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05134_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] _00846_ vssd1 vssd1
+ vccd1 vccd1 _00847_ sky130_fd_sc_hd__xnor2_1
Xhold424 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\] vssd1 vssd1
+ vccd1 vccd1 net1094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\] vssd1 vssd1
+ vccd1 vccd1 net1105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\] vssd1 vssd1 vccd1
+ vccd1 net1127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 team_07_WB.instance_to_wrap.team_07.label_num_bus\[3\] vssd1 vssd1 vccd1
+ vccd1 net1138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05065_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up vssd1 vssd1
+ vccd1 vccd1 _00794_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09942_ net463 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
Xhold479 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[0\] _04870_ vssd1
+ vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06529__A2 _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _04141_ _04170_ net196 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__a21oi_1
X_08755_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[29\] net1158 net236 vssd1
+ vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__mux2_1
X_05967_ net260 net214 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__nor2_1
X_07706_ _01735_ _01901_ net188 vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__o21a_1
X_04918_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
X_08686_ net1152 _04105_ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__a21oi_1
X_05898_ _01565_ _01569_ _01570_ _01573_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__or4_1
X_07637_ _03152_ _03178_ _03194_ _03099_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07568_ _02150_ _02191_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09307_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[10\]
+ _04491_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__or2_1
X_06519_ _02153_ _02189_ _02190_ _02192_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_63_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07499_ net93 _02348_ _02343_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09238_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__inv_2
XANTENNA__07500__B _02673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05301__A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04391_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06116__B net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06217__A1 _01600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05020__B net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08612__A _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06768__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05955__B net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07178__C1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07717__A1 _01649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ clknet_leaf_42_wb_clk_i _00092_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08758__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05971__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05690__B _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10915_ net660 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_98_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10846_ net522 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10777_ clknet_leaf_65_wb_clk_i _00598_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07545__A1_N _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05211__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07956__A1 _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05865__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06042__A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07708__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10560__Q team_07_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05982__A3 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06870_ _02535_ _02540_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05821_ _01494_ _01497_ _01514_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08540_ _03628_ _03650_ net146 vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09072__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05752_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\] _01450_ vssd1 vssd1
+ vccd1 vccd1 _01451_ sky130_fd_sc_hd__or4b_1
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08471_ net486 net488 _03710_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__or3b_1
X_05683_ net441 net440 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_46_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07422_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\]
+ _03004_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07353_ _00708_ _00816_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10753__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06304_ net199 _01977_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_135_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07284_ _02917_ _02918_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[10\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_135_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09023_ net251 _04282_ _04284_ net405 net994 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06235_ net91 _01670_ _01706_ _01912_ _01913_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__o32a_1
XFILLER_0_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout307_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold210 _00500_ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__dlygate4sd3_1
X_06166_ _01832_ _01836_ _01838_ _01846_ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__a211o_1
Xhold221 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold232 team_07_WB.instance_to_wrap.team_07.label_num_bus\[33\] vssd1 vssd1 vccd1
+ vccd1 net902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold243 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__dlygate4sd3_1
X_05117_ _00685_ _00828_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__and2_1
Xhold254 _00474_ vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__dlygate4sd3_1
X_06097_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[14\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\]
+ _01779_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__or3_1
Xhold265 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\] vssd1 vssd1
+ vccd1 vccd1 net935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06223__Y _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold276 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[5\] vssd1 vssd1
+ vccd1 vccd1 net946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold287 _00093_ vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__dlygate4sd3_1
X_05048_ _00768_ _00769_ _00770_ _00779_ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09925_ net935 _01784_ _04870_ _04902_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__o31ai_1
Xhold298 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[20\]
+ vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09856_ _04827_ _04859_ vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__nor2_1
X_08807_ net195 _04159_ vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__nor2_1
XANTENNA__05186__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06383__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09787_ _00657_ _04803_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__nor2_2
X_06999_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\] _02654_
+ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__xor2_1
X_10985__626 vssd1 vssd1 vccd1 vccd1 _10985__626/HI net626 sky130_fd_sc_hd__conb_1
X_08738_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__mux2_1
XANTENNA__07537__D_N _03095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ _04080_ _04095_ _04084_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__o21ai_1
X_10700_ clknet_leaf_69_wb_clk_i _00531_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05015__B net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10631_ clknet_leaf_50_wb_clk_i _00495_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09624__A1 _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10562_ clknet_leaf_24_wb_clk_i _00430_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06127__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10493_ clknet_leaf_15_wb_clk_i _00361_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05966__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09927__A2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06414__X _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06374__B1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06126__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06677__A1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10829_ net505 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_138_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06429__A1 _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06020_ net106 net142 net169 net205 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07929__A1 _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07929__B2 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08051__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06601__A1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07971_ _03377_ _03405_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__nor2_1
X_09710_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\] _04752_ vssd1
+ vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__and2_1
X_06922_ _02591_ _02592_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__or2_1
XANTENNA__09551__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__or4b_1
X_06853_ _02499_ _02504_ _02507_ net190 _02523_ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__o221a_1
XANTENNA__05168__B2 team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05804_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\] _01486_
+ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__nand2_1
X_09572_ net480 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _04657_ _04660_ vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06784_ _02431_ _02454_ _02455_ _02428_ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08523_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\]
+ _03983_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__and3_1
X_05735_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\] _00787_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout257_A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ _03667_ _03826_ _03923_ _03926_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06668__B2 _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04955__A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05666_ net419 _00676_ _00677_ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_137_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07405_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] _02994_
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[8\] vssd1 vssd1 vccd1
+ vccd1 _02997_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_102_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08385_ _03718_ _03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout424_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05597_ _01302_ _01303_ _01304_ _01309_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07336_ _02414_ _02948_ _01175_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07267_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09006_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06218_ _01894_ _01895_ _01897_ _01889_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07198_ _02773_ _02846_ _02781_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06149_ net102 _01828_ net214 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05946__A3 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ net1103 net154 net152 _04892_ vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__a22o_1
XANTENNA__07148__A2 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ _04824_ _04845_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_126_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07608__B1 _01672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10614_ clknet_leaf_54_wb_clk_i _00478_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08771__S net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07084__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10545_ clknet_leaf_18_wb_clk_i _00413_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10476_ clknet_leaf_17_wb_clk_i _00344_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08336__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06347__B1 _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06898__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05520_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ _01219_ _01232_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_129_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05322__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05451_ _01042_ _01068_ _01102_ _01020_ vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_16 team_07_WB.instance_to_wrap.team_07.recFLAG.flagDetect vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_27 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ net466 _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05382_ _00970_ _01063_ vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07121_ _01635_ _02757_ _02769_ _02774_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07052_ _02677_ _02691_ _02706_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06003_ net219 net198 _01682_ _01695_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__o31a_2
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07954_ _01057_ _01658_ _03369_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__a21o_1
XANTENNA__08327__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06905_ net433 net182 net173 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__o2bb2a_1
X_07885_ net267 _03285_ _03413_ _03439_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout374_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ _04666_ _04692_ _04693_ _04664_ net1071 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__a32o_1
X_06836_ net432 _02506_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__nor2_1
XANTENNA__05010__A0 team_07_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07550__A2 _02262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09555_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[47\]
+ net225 _04605_ net887 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_06767_ net280 net430 net278 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_104_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout162_X net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\]
+ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__and3_1
X_05718_ net483 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[16\]
+ net270 _04617_ net291 net223 vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06698_ net177 _02274_ net258 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_121_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08437_ _00711_ _00727_ _03717_ _03910_ _00048_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_93_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05649_ _01360_ _01361_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07996__A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08368_ _00729_ _01380_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09055__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07319_ _01190_ _01192_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08299_ net5 _00663_ _03703_ _03705_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a41o_2
XFILLER_0_6_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05077__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10330_ clknet_leaf_52_wb_clk_i net688 net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_10261_ clknet_leaf_74_wb_clk_i _00253_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10192_ clknet_leaf_84_wb_clk_i _00196_ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05963__B net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout350 net389 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_128_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout361 net363 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07236__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout372 net374 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06329__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout383 net384 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_2
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout394 _03562_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__buf_2
XFILLER_0_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__B1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05978__X _01672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05855__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07057__A1 _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09987__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput36 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
X_10528_ clknet_leaf_25_wb_clk_i _00396_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06804__B2 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ clknet_leaf_22_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_left
+ net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06034__B _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06050__A _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04951_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07670_ net104 _02277_ _03173_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__o21a_1
X_06621_ _01698_ _02021_ net258 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__o21ai_4
XANTENNA__10344__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09340_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__a31o_1
X_06552_ _01618_ net253 _02196_ net265 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05503_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ _01215_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__xnor2_1
X_09271_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ _04467_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__or3b_1
X_06483_ _02155_ _02156_ _02153_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08222_ team_07_WB.instance_to_wrap.team_07.buttonHighlightPixel _00728_ team_07_WB.instance_to_wrap.team_07.buttonPixel
+ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05434_ _00982_ _01027_ _01091_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08153_ net471 _00717_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05365_ net397 _01056_ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__nand2_4
XFILLER_0_126_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout122_A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07104_ net82 _02756_ _02757_ _01635_ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__o211a_4
XFILLER_0_28_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05400__Y _01113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08084_ net898 _03594_ _03595_ net956 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05296_ _01001_ _01008_ vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__or2_1
XANTENNA__06225__A _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10161__RESET_B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07035_ _02688_ _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_77_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout491_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06023__A2 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ _04255_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__or4_1
X_07937_ _03487_ _03491_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07868_ net397 _01058_ _02106_ _00749_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_3_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07523__A2 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09607_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[10\]
+ _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06819_ net111 _02477_ _02478_ _02488_ _02489_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__o221a_1
XANTENNA__05534__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07799_ _03340_ _03346_ _03353_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__or3_2
XFILLER_0_35_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09538_ net291 _04645_ _04649_ net271 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[36\]
+ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05638__A_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09469_ net928 net207 _04607_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05023__B net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07039__A1 _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05958__B net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08236__B1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06406__Y _02080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ clknet_leaf_45_wb_clk_i net759 net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_11019__643 vssd1 vssd1 vccd1 vccd1 _11019__643/HI net643 sky130_fd_sc_hd__conb_1
XFILLER_0_81_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05974__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05470__B1 _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ clknet_leaf_82_wb_clk_i _00236_ net319 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07211__A1 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10175_ clknet_leaf_8_wb_clk_i _00185_ net329 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06905__A2_N net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850__526 vssd1 vssd1 vccd1 vccd1 _10850__526/HI net526 sky130_fd_sc_hd__conb_1
XANTENNA__07762__A2 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout180 _01544_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_4
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07514__A2 _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05525__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08475__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05150_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[2\] _00862_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__mux2_4
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05081_ net412 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ sky130_fd_sc_hd__inv_6
XANTENNA__05461__B1 _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _04143_ _04180_ _04144_ vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07202__B2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06051__Y _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08771_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[5\] net713 net245 vssd1
+ vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__mux2_1
X_05983_ net163 net149 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__nor2_4
XANTENNA__06961__B1 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ _01064_ net115 vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__nor2_1
X_04934_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07604__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ _03063_ _03064_ _03210_ _03209_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__o31a_1
X_06604_ _01651_ _01936_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__nor2_4
XFILLER_0_88_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07584_ _02232_ _03142_ _02830_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_76_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09323_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ _04502_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06535_ net268 net276 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout337_A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09254_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ _04454_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07674__D1 _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06466_ net277 _02030_ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_32_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08205_ net421 team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] _01258_
+ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05417_ _00668_ _01055_ _01129_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__a21oi_1
X_09185_ _04404_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__inv_2
X_06397_ net166 _02069_ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout125_X net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[21\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[20\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\]
+ _03621_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__or4_2
X_05348_ net194 _01000_ _01004_ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__or3_2
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08067_ net456 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05279_ _00979_ _00987_ vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07018_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[2\] _00828_ vssd1 vssd1
+ vccd1 vccd1 _02673_ sky130_fd_sc_hd__nor2_2
XFILLER_0_113_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08170__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10953__594 vssd1 vssd1 vccd1 vccd1 _10953__594/HI net594 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_52_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08969_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\] net782
+ net448 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05018__B net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ net581 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_116_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10862_ net538 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10793_ clknet_leaf_75_wb_clk_i _00614_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05969__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10083__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07680__A1 net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10012__RESET_B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05443__B1 _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05994__A1 _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891__648 vssd1 vssd1 vccd1 vccd1 net648 _10891__648/LO sky130_fd_sc_hd__conb_1
X_10227_ clknet_leaf_0_wb_clk_i _00231_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09463__X _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05991__X _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ clknet_leaf_2_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[5\]
+ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[3\]
+ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__dlygate4sd3_1
X_10089_ clknet_leaf_68_wb_clk_i _00147_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07499__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06320_ net177 _01973_ _01984_ _01986_ _01976_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a41o_1
XFILLER_0_127_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06251_ _01927_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07671__A1 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07671__B2 _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06046__Y _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05202_ _00907_ _00914_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06182_ _01858_ _01860_ _01861_ _01862_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_96_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold403 team_07_WB.instance_to_wrap.team_07.label_num_bus\[7\] vssd1 vssd1 vccd1
+ vccd1 net1073 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold414 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__dlygate4sd3_1
X_05133_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[8\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\]
+ _00843_ _00840_ vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__mux4_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold425 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold436 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\] vssd1 vssd1
+ vccd1 vccd1 net1106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold447 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold458 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold469 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[4\] vssd1 vssd1
+ vccd1 vccd1 net1139 sky130_fd_sc_hd__dlygate4sd3_1
X_05064_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right vssd1
+ vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09941_ net463 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06503__A _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ net341 _01790_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_111_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08823_ net831 _04169_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__nand2_1
XANTENNA__06934__B1 _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout287_A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08754_ net1143 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__mux2_1
X_05966_ net260 _01659_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__nor2_4
X_07705_ net167 net103 vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__nand2_1
X_04917_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] vssd1 vssd1
+ vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
X_08685_ _04049_ _04073_ _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__and3_1
X_05897_ _01562_ net147 _01572_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout454_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07636_ _02061_ _03193_ _03165_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06162__A1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06162__B2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07567_ _02217_ _02223_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__nor2_1
X_09306_ net229 _04490_ _04492_ net404 net1125 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06518_ _02108_ _02150_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07498_ _00943_ _02250_ _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__and3b_1
XFILLER_0_134_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09237_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04418_ _04435_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_118_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06449_ _01686_ _01703_ _01722_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09168_ net210 _04390_ _04392_ net401 net807 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08119_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[1\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[0\] vssd1
+ vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__or2_1
XANTENNA__06116__C _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05795__Y _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09099_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04318_ _04333_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05425__B1 _01113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08104__S _02671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07178__B1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ clknet_leaf_58_wb_clk_i _00009_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05728__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05971__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input15_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10914_ net659 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XANTENNA__08774__S net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06153__A1 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10845_ net521 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10776_ clknet_leaf_65_wb_clk_i _00597_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08850__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07956__A2 _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10856__532 vssd1 vssd1 vccd1 vccd1 _10856__532/HI net532 sky130_fd_sc_hd__conb_1
XFILLER_0_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06042__B _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05820_ _01495_ _01496_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05751_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\] _01449_ vssd1 vssd1
+ vccd1 vccd1 _01450_ sky130_fd_sc_hd__nor4_1
XFILLER_0_77_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08470_ _00729_ _03940_ _03941_ _03738_ net486 vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__a311o_1
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05682_ _01318_ _01393_ _01394_ vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__nand3_1
X_07421_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\]
+ _03003_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\] vssd1
+ vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07352_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[18\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[16\] _02958_
+ _02960_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_98_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06303_ net216 _01967_ _01968_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__or3_1
XANTENNA__05402__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07283_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_135_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09022_ _04283_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06234_ net114 _01880_ _01911_ net91 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold200 _00484_ vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06165_ _01839_ _01845_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout202_A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold222 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[24\] vssd1 vssd1
+ vccd1 vccd1 net892 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06504__Y _02178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold233 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[7\]
+ vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__dlygate4sd3_1
X_05116_ _00685_ _00828_ vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__nor2_2
Xhold244 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[27\]
+ vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[37\]
+ vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__dlygate4sd3_1
X_06096_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[12\] _01778_
+ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold266 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[17\]
+ vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[45\]
+ vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold288 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[20\] vssd1 vssd1
+ vccd1 vccd1 net958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\] vssd1 vssd1
+ vccd1 vccd1 net969 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _01784_ net155 net935 vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__o21ai_1
X_05047_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[8\]
+ _00777_ _00778_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input7_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ net247 _04858_ _04857_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06520__X _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10775__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ net1060 _04158_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__xnor2_1
X_06998_ _02655_ _02656_ _02661_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__and3_1
XANTENNA__06383__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09786_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__nand2_1
XANTENNA__07064__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08737_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ net234 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__mux2_1
X_05949_ net214 _01642_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__nand2_1
X_08668_ _04089_ _04092_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__and2b_1
XANTENNA__07332__A0 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07619_ net254 _01731_ _02271_ _03114_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08599_ _03624_ _04033_ net146 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06150__A4 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10630_ clknet_leaf_49_wb_clk_i _00494_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06408__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10561_ clknet_leaf_24_wb_clk_i _00429_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07635__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08832__B1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06127__B _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10492_ clknet_leaf_15_wb_clk_i _00360_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06143__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08769__S net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06374__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__B1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10445__RESET_B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06677__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10927__577 vssd1 vssd1 vccd1 vccd1 _10927__577/HI net577 sky130_fd_sc_hd__conb_1
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10828_ net504 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06429__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10759_ clknet_leaf_67_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[6\]
+ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10897__654 vssd1 vssd1 vccd1 vccd1 net654 _10897__654/LO sky130_fd_sc_hd__conb_1
XFILLER_0_23_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07929__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08051__A1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06053__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06601__A2 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ _01692_ _03385_ _03524_ _03523_ _01651_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__o32a_1
XANTENNA__08055__A_N net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06921_ net432 net182 _02509_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__and3_1
X_09640_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _04702_ _00761_
+ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__o21ai_1
X_06852_ net432 net182 _02506_ _02517_ _02522_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__o311a_1
X_05803_ _01495_ _01496_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__and2_1
X_09571_ _04657_ _04625_ _04612_ _01421_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__and4b_1
X_06783_ _02426_ _02450_ _02451_ _02448_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__o2bb2a_1
X_08522_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\] _03983_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05734_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\] _01437_ _01438_
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[0\]
+ sky130_fd_sc_hd__a21bo_1
XANTENNA__08708__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ _03925_ _03630_ _03631_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_65_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05665_ _01371_ _01377_ net442 _01322_ _01370_ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_137_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07404_ net1000 _02994_ _02996_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[7\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08384_ _03739_ _03805_ _03723_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_82_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05596_ _01303_ _01304_ _01307_ _01308_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_102_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05132__A team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07617__A1 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07335_ _02413_ _02947_ _00965_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07266_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09005_ _04253_ net251 _04271_ net403 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06217_ _01600_ _01824_ _01896_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__o21bai_1
X_07197_ _02040_ _02775_ _02836_ _02848_ _02767_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__a32o_1
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout205_X net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07059__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06148_ net176 _01723_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__nand2_2
X_06079_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\] _01763_ _01764_
+ _01765_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__and4_1
X_09907_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\] _01779_
+ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__xnor2_1
X_09838_ net269 _04845_ _04846_ net247 net1048 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09769_ _04794_ _04795_ vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_126_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05026__B _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07856__B2 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06513__D1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07608__A1 _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10613_ clknet_leaf_49_wb_clk_i _00477_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10544_ clknet_leaf_18_wb_clk_i _00412_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07084__A2 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10475_ clknet_leaf_17_wb_clk_i _00343_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06044__B1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10697__RESET_B net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05983__Y _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output46_A net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07847__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05450_ _01009_ _01076_ _01103_ _01069_ vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__o22a_1
XANTENNA__08962__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06048__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_28 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05381_ net299 _01062_ vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__nor2_4
XFILLER_0_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07120_ net88 _02109_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07051_ _01902_ _02087_ _02695_ _02705_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a31o_1
XFILLER_0_125_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06002_ net170 net104 _01693_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06511__A _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ net277 _03355_ _03356_ _03506_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__or4_1
XFILLER_0_103_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06904_ _02534_ _02574_ _02532_ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a21oi_1
X_07884_ _03285_ _03438_ _03282_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_108_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09623_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\]
+ _04688_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__nand3_1
X_06835_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout367_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ net887 net209 _04656_ vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__o21a_1
X_06766_ net90 _02413_ _02437_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_104_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07342__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__nor4_1
XFILLER_0_66_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05717_ _01412_ _01413_ _01425_ _01428_ net246 vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_19_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06697_ _02214_ _02258_ _02362_ net265 _02190_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a221o_1
X_09485_ _04613_ _04616_ _00667_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_121_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08436_ _03835_ _03909_ net489 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__a21o_1
X_05648_ _00678_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] _01359_ vssd1
+ vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_77_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08872__S net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08367_ net459 _01270_ _01296_ _01302_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wireHighlightPixel
+ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__a41o_1
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05579_ _01281_ _01289_ _01290_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07318_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[1\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08298_ net416 _03775_ net488 vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05077__B2 _00675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07249_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06405__B net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10260_ clknet_leaf_74_wb_clk_i _00252_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06124__C _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10191_ clknet_leaf_90_wb_clk_i _00195_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06577__A1 _02178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07517__A _03075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout340 net341 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout351 net357 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_4
Xfanout362 net363 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07236__B _02082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout373 net374 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_2
XANTENNA__06329__A1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout384 net388 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout395 net396 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_2
XFILLER_0_69_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07829__A1 _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07829__B2 _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput15 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07057__A2 _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput26 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput37 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10527_ clknet_leaf_21_wb_clk_i _00395_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09203__A0 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10458_ clknet_leaf_22_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.edge_back
+ net338 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_21_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06568__A1 _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10389_ clknet_leaf_11_wb_clk_i net770 net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04950_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_53_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06050__B _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__S _04245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06620_ _02280_ _02292_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06551_ _02220_ _02222_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_48_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05502_ net422 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_75_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09270_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04420_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__or4b_1
XANTENNA__10639__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06482_ net103 _02056_ _02054_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08221_ team_07_WB.instance_to_wrap.team_07.heartPixel team_07_WB.instance_to_wrap.team_07.labelPixel\[1\]
+ _03699_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__or3_4
X_05433_ _01059_ _01060_ _01144_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05888__Y _01582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08152_ net473 _03635_ _03637_ _03634_ vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05364_ net437 _01049_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06506__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07103_ _02249_ net82 vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08083_ net956 net232 _03595_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__a22o_1
X_05295_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[2\]
+ net427 _00988_ _00980_ vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_28_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout115_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06225__B _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07034_ _02085_ _02185_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06241__A _01672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__or4b_1
X_07936_ net256 _03475_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ net274 _03392_ _03395_ _03396_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__or4_1
XANTENNA__04967__Y _00706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09606_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\]
+ _04675_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_123_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06818_ _02478_ _02488_ net118 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__a21o_1
XANTENNA__08168__A _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07798_ _03347_ _03350_ _03351_ _03352_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__or4_1
XFILLER_0_74_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09537_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\] _01420_
+ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__or2_1
X_06749_ _00672_ net150 net159 net428 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09468_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[9\]
+ net273 net292 net222 vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07800__A _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08419_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\] _00704_
+ _03646_ _03893_ _03630_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a41o_1
X_09399_ _04556_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08236__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06135__B _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10312_ clknet_leaf_45_wb_clk_i net737 net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_15_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10243_ clknet_leaf_86_wb_clk_i _00235_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__05974__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ clknet_leaf_9_wb_clk_i _00184_ net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06151__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout170 _01685_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_4
Xfanout181 _01643_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_4
Xfanout192 _01003_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_2
XANTENNA__06707__D1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06486__B1 _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07683__C1 _01905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08227__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05080_ team_07_WB.EN_VAL_REG _00065_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10311__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[4\] net878 net245 vssd1
+ vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__mux2_1
X_05982_ net156 net131 net124 net137 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__a31o_4
XTAP_TAPCELL_ROW_72_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07721_ _03274_ _03275_ _03273_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__o21bai_2
X_04933_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07604__B _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ _01904_ _02278_ _03188_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__o21a_1
XANTENNA__06713__A1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06603_ _02275_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__inv_2
X_07583_ _01655_ _01717_ _01828_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09322_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[14\]
+ _04502_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06534_ _02129_ _02150_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09253_ net230 _04453_ _04455_ net406 net950 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06465_ net277 _02030_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__nor2_2
XFILLER_0_75_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08204_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\]
+ _00730_ _01260_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__and4_1
X_05416_ _00966_ _01089_ _01128_ _01064_ _01075_ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09184_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ _04399_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06396_ _01676_ _01688_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08135_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\]
+ _03621_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_79_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05347_ _01000_ net191 _01021_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout118_X net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ net395 net296 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ _03586_ vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_116_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05278_ net193 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07017_ net943 _02672_ _02670_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10873__549 vssd1 vssd1 vccd1 vccd1 _10873__549/HI net549 sky130_fd_sc_hd__conb_1
X_08968_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[8\] net810
+ net448 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__mux2_1
X_07919_ _03305_ _03445_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__nor2_1
X_08899_ net481 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[6\] vssd1
+ vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__and3_1
X_10930_ net580 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__07901__B1 _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10861_ net537 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_67_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06180__A2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10792_ clknet_leaf_77_wb_clk_i _00613_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05969__B _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07680__A2 _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05985__A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10226_ clknet_leaf_85_wb_clk_i _00230_ net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\]
+ sky130_fd_sc_hd__dfrtp_4
X_10157_ clknet_leaf_2_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[4\]
+ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06943__A1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[8\]
+ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_50_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07705__A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10088_ clknet_leaf_66_wb_clk_i _00146_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07499__A2 _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_X clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06250_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] net458 vssd1 vssd1
+ vccd1 vccd1 _01927_ sky130_fd_sc_hd__nand2_1
XANTENNA__08970__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05201_ _00912_ _00913_ _00911_ vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__or3b_1
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06181_ _00649_ net133 net121 _00635_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_96_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05132_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] _00844_ vssd1 vssd1
+ vccd1 vccd1 _00845_ sky130_fd_sc_hd__xnor2_1
Xhold404 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold415 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[34\]
+ vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 team_07_WB.instance_to_wrap.team_07.label_num_bus\[4\] vssd1 vssd1 vccd1
+ vccd1 net1096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold437 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[2\] vssd1 vssd1
+ vccd1 vccd1 net1107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold448 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] vssd1 vssd1
+ vccd1 vccd1 net1118 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05063_ _00792_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[2\]
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_74_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09940_ net463 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
Xhold459 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06503__B _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09871_ net411 _01789_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07187__A1 _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _04168_ _04169_ net196 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07615__A _02873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08753_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[27\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ net235 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__mux2_1
X_05965_ net214 _01656_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout182_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07704_ _01683_ _02046_ _03259_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__or3_1
X_04916_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _00656_ sky130_fd_sc_hd__inv_2
X_08684_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared _04081_ vssd1
+ vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__nor2_1
X_05896_ _01585_ _01589_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__nand2_2
XANTENNA__09884__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06698__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ net135 _01683_ _01687_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout447_A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07566_ _03106_ _03116_ _03119_ _03124_ _03104_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__a221o_1
XANTENNA__05370__B1 _01067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09305_ _04491_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07647__C1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06517_ net282 _02106_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__and2_4
XFILLER_0_119_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07497_ _01640_ _03053_ _03056_ _02390_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__a2bb2o_1
X_09236_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[7\]
+ _04440_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_118_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06448_ _01693_ _02047_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09167_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06379_ _01687_ _01690_ _01696_ _02052_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__o31a_1
XFILLER_0_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08118_ net832 net814 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09098_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04333_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[19\]
+ net394 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout95_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07178__A1 _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ clknet_leaf_55_wb_clk_i _00008_ net360 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05728__A2 _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07525__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10913_ net658 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06153__A2 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10844_ net520 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05699__B _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10775_ clknet_leaf_65_wb_clk_i _00596_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06147__Y _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08643__X _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05986__Y _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06604__A _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05416__B2 _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10209_ clknet_leaf_81_wb_clk_i _00213_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08030__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05750_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[5\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__or4_1
XANTENNA__08965__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09330__A2 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05681_ net441 _01392_ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07420_ net1050 _03004_ _03006_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[13\]
+ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07351_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[20\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[19\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06302_ _01967_ _01968_ net216 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05402__B _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07282_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ _00679_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09021_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ _04280_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__and2_1
X_06233_ _01865_ _01870_ _01880_ _01614_ _01882_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_135_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06164_ _01820_ _01842_ _01844_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a21oi_1
Xhold201 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06073__X _01760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold212 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold223 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[6\]
+ vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05115_ team_07_WB.instance_to_wrap.team_07.memGen.stage\[1\] net450 vssd1 vssd1
+ vccd1 vccd1 _00828_ sky130_fd_sc_hd__or2_2
XFILLER_0_41_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold234 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[18\]
+ vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__dlygate4sd3_1
X_06095_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[11\]
+ _01777_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__or3_1
XANTENNA__08947__A_N net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold245 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[11\]
+ vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold256 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[21\]
+ vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold267 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[35\]
+ vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[36\]
+ vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _01784_ _04870_ _04901_ vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__o21ai_1
X_05046_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\] vssd1 vssd1 vccd1 vccd1
+ _00778_ sky130_fd_sc_hd__or3b_1
XFILLER_0_102_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold289 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[5\] vssd1 vssd1
+ vccd1 vccd1 net959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09854_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[14\] _04855_ vssd1
+ vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__nand2_1
X_08805_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[8\] _04156_ vssd1
+ vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__nor2_1
X_09785_ _00657_ _04809_ _04808_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__a2bb2o_1
X_06997_ _02658_ _02660_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__or2_1
XANTENNA__06383__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout185_X net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ net238 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__mux2_1
XANTENNA__07064__B _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05948_ net260 net197 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__nor2_2
XFILLER_0_96_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08667_ _04076_ _04094_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05879_ _01562_ net147 _01564_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07618_ _02208_ _03127_ _03128_ _03175_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__o31a_1
X_08598_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ _03623_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07080__A _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05894__A1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ _02838_ _03107_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05312__B _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10560_ clknet_leaf_89_wb_clk_i _00428_ _00065_ vssd1 vssd1 vccd1 vccd1 team_07_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07635__A2 _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10922__667 vssd1 vssd1 vccd1 vccd1 net667 _10922__667/LO sky130_fd_sc_hd__conb_1
XANTENNA__06127__C _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ _04430_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10491_ clknet_leaf_15_wb_clk_i _00359_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__A1_N net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10879__555 vssd1 vssd1 vccd1 vccd1 _10879__555/HI net555 sky130_fd_sc_hd__conb_1
XFILLER_0_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout98_X net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07571__A1 _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06374__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06126__A2 _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07874__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05885__A1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10827_ net503 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_7_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05997__X _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10758_ clknet_leaf_61_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[5\]
+ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06605__Y _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10689_ clknet_leaf_53_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[21\]
+ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06053__B net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06920_ net174 _02511_ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09551__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ _02521_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05802_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\]
+ _01486_ _01487_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__and4_2
X_09570_ net480 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ _04657_ _04659_ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_69_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06782_ net428 net159 _02445_ _02453_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08521_ net873 _03982_ vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05733_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\] _00772_ _00784_
+ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__or3_1
XFILLER_0_136_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08452_ _03924_ _03892_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_65_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05664_ _01256_ _01259_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_137_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07403_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\] _02994_
+ net478 vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09067__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ net490 _03855_ _03858_ _03751_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__o31a_1
X_05595_ net420 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] vssd1 vssd1 vccd1
+ vccd1 _01308_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_102_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout145_A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07334_ net430 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__mux2_1
XANTENNA__07617__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05628__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07265_ _02905_ _02906_ _01315_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[15\]
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout312_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09004_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06216_ _01850_ _01893_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__nand2_1
X_07196_ net160 _01688_ _02836_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06244__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06147_ net173 _01724_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__nor2_4
XANTENNA__07059__B _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10991__632 vssd1 vssd1 vccd1 vccd1 _10991__632/HI net632 sky130_fd_sc_hd__conb_1
X_06078_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\] vssd1 vssd1 vccd1
+ vccd1 _01765_ sky130_fd_sc_hd__nor3_1
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09906_ net848 net154 net152 _04891_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__a22o_1
X_05029_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05147__X _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ _04838_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\] vssd1 vssd1
+ vccd1 vccd1 _04846_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07553__A1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05307__B _01014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ _04767_ _04790_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ net962 _04132_ _04133_ vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__a21oi_1
X_09699_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\] net250 _04742_
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\] vssd1 vssd1 vccd1
+ vccd1 _04747_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07522__B _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06513__C1 _01660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10612_ clknet_leaf_49_wb_clk_i _00476_ net371 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07608__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10543_ clknet_leaf_18_wb_clk_i _00411_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05977__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07084__A3 _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06425__Y _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10474_ clknet_leaf_14_wb_clk_i _00342_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06044__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05993__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07544__A1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10666__RESET_B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05217__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06048__B _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05380_ _01002_ _01023_ _01092_ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__o21ai_1
XANTENNA_18 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_29 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05887__B _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07050_ _02692_ _02701_ _02704_ _02699_ _02703_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a221o_1
XANTENNA__06283__A1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10975__616 vssd1 vssd1 vccd1 vccd1 _10975__616/HI net616 sky130_fd_sc_hd__conb_1
X_06001_ net133 net121 _01676_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06035__A1 _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06860__A1_N net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07952_ net274 _03346_ _03506_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__or3b_1
XANTENNA__06511__B _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06903_ _02538_ _02573_ _02536_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__o21bai_1
X_07883_ _02331_ _03291_ _03290_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_108_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09622_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\] _04688_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_108_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06834_ _02504_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09553_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[45\]
+ net273 net293 net224 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a211o_1
X_06765_ _02430_ _02435_ _02436_ _02426_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout262_A _01488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08504_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\]
+ _00697_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[11\] vssd1 vssd1
+ vccd1 vccd1 _03970_ sky130_fd_sc_hd__and4b_1
XFILLER_0_37_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05716_ net414 _01411_ _01423_ _00826_ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__and4bb_1
X_09484_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] vssd1
+ vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__nand2b_1
X_06696_ _02271_ _02364_ _02365_ _02367_ _02368_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a32o_1
XANTENNA__06239__A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08435_ net486 _03846_ _03873_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__or3_1
X_05647_ _00678_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\] _01359_ vssd1
+ vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_121_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout148_X net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08366_ _01253_ _01381_ _03733_ _03841_ net460 vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__o32a_1
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05578_ _01289_ _01290_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__and2_1
XANTENNA__08799__B1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07317_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ _00723_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_y\[2\]
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_18_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08297_ net459 _03774_ _03694_ _00729_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07248_ _02893_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[4\]
+ _02895_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[4\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_46_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06405__C _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07179_ _02822_ _02826_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__or2_1
X_10190_ clknet_leaf_84_wb_clk_i _00194_ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06702__A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__B2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout330 net339 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_4
Xfanout341 net389 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_128_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout352 net357 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_4
Xfanout363 net388 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__clkbuf_4
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_2
Xfanout385 net387 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__clkbuf_4
Xfanout396 _03024_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07533__A _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07829__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05988__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06436__X _02110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_5_0_wb_clk_i_X clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput16 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput27 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06265__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10526_ clknet_leaf_21_wb_clk_i _00394_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10457_ clknet_leaf_13_wb_clk_i _00337_ net335 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08652__B1_N _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10388_ clknet_leaf_11_wb_clk_i net696 net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_103_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06568__A2 _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08962__A0 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11009_ net639 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06550_ _01611_ net253 _02223_ _02043_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__or4b_1
XANTENNA__08973__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05501_ net422 _00691_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ _01198_ _01213_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_16_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06481_ _01828_ _02154_ net203 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08220_ team_07_WB.instance_to_wrap.team_07.labelPixel\[0\] team_07_WB.instance_to_wrap.team_07.labelPixel\[3\]
+ team_07_WB.instance_to_wrap.team_07.labelPixel\[2\] team_07_WB.instance_to_wrap.team_07.displayPixel
+ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05432_ _01144_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
XANTENNA__06346__X _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08274__A net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003__638 vssd1 vssd1 vccd1 vccd1 _11003__638/HI net638 sky130_fd_sc_hd__conb_1
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08151_ _00717_ net472 vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__nor2_2
X_05363_ net437 _01049_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__nor2_2
XANTENNA__06506__B net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07102_ net265 _02197_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07453__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08082_ net482 _00815_ _03593_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__and3_2
X_05294_ _01002_ _01006_ vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07033_ _01636_ net83 _02350_ _02335_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout108_A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06522__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06559__A2 _02230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10588__RESET_B net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08984_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[13\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ _04253_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__or3_1
X_07935_ _03479_ _03488_ _03489_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__and3b_1
XANTENNA__07508__A1 _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08705__B1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07866_ _03339_ _03419_ _03420_ _03397_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09605_ _03976_ _04679_ _04680_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_123_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06817_ net274 _02487_ _02482_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_123_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07797_ _01115_ net111 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout265_X net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ net948 net206 _04648_ vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06748_ net174 _02418_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ net945 net208 _04606_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06679_ _00759_ net84 _02250_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08418_ _03655_ _03891_ _03892_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07800__B net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ net414 _04555_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__or2_2
XANTENNA__06523__C_N _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08349_ net470 _03660_ net467 vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_19_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08236__A2 _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08912__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10311_ clknet_leaf_45_wb_clk_i net733 net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_120_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10242_ clknet_leaf_86_wb_clk_i _00234_ net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06432__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10173_ clknet_leaf_9_wb_clk_i _00183_ net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input38_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 _01557_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_8
Xfanout171 _01681_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_4
Xfanout182 net183 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_4
Xfanout193 net194 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08172__B2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08646__X _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08381__X _03857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10509_ clknet_leaf_16_wb_clk_i _00377_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08033__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08968__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05981_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[1\] _01633_ vssd1
+ vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_72_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08950__A3 _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06961__A2 _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ _01105_ _01597_ _01604_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__and3_1
X_04932_ net429 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07651_ _03098_ _03099_ _03207_ _03208_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__a22o_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07604__C _03162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06174__B1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07910__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06602_ net175 _02013_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__nand2_1
X_07582_ _02842_ _03140_ _03118_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09321_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[13\]
+ _04499_ _04501_ _04503_ vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__o22a_1
XANTENNA__10756__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06533_ _02102_ _02155_ _02153_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__inv_2
X_06464_ net278 net277 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__nor2_2
XFILLER_0_47_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06517__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08203_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\] _00730_ vssd1
+ vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05415_ _01023_ _01100_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__nor2_1
X_09183_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[10\]
+ _04396_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_32_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06395_ _01677_ _01689_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout225_A _04582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08134_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[18\]
+ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__or2_1
X_05346_ net193 _01000_ _01019_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_79_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08065_ net453 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05277_ _00982_ _00988_ _00989_ vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_116_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07016_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\]
+ _02671_ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08967_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[7\] net816
+ net448 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__mux2_1
X_07918_ _01083_ net147 _03443_ _03441_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__a31o_1
X_08898_ _04214_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[6\]
+ _04209_ vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__mux2_1
XANTENNA__09351__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07849_ _00747_ _03354_ _03363_ net268 vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__o22a_1
XANTENNA__07901__A1 _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ net536 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_66_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09519_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[31\]
+ net222 _04605_ net896 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07811__A _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10791_ clknet_leaf_77_wb_clk_i _00612_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06468__A1 _02119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06468__B2 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_61_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06427__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09964__SET_B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07680__A3 _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07968__A1 _01113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08090__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05985__B net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05979__B1 _01672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06433__Y _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10225_ clknet_leaf_0_wb_clk_i _00229_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10156_ clknet_leaf_2_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[3\]
+ net309 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold5 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07705__B net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ clknet_leaf_69_wb_clk_i _00145_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload3_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10989_ net630 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_48_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05593__C_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05200_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] _00901_ vssd1 vssd1
+ vccd1 vccd1 _00913_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06180_ net289 net136 _01859_ _01860_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_96_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05131_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[9\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\]
+ _00843_ _00840_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__mux4_2
Xhold405 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\] vssd1 vssd1
+ vccd1 vccd1 net1075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold427 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\] vssd1
+ vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07168__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold438 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[8\] vssd1 vssd1 vccd1
+ vccd1 net1108 sky130_fd_sc_hd__dlygate4sd3_1
X_05062_ _00785_ _00789_ _00790_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__nand3_1
Xhold449 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\] vssd1 vssd1
+ vccd1 vccd1 net1119 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06072__A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08908__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09870_ _00827_ _01789_ net411 vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[14\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\]
+ _01448_ _04160_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_5_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06934__A2 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08752_ net1157 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__mux2_1
X_05964_ _01503_ net197 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__nand2_4
X_07703_ _01686_ _01737_ _02040_ _01646_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04915_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _00655_ sky130_fd_sc_hd__inv_2
X_08683_ _04106_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ _04105_ vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__mux2_1
X_05895_ _01586_ _01588_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout175_A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07634_ net103 _02056_ _02085_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__o21ba_1
XANTENNA__06698__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06162__A3 _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ _01704_ _02219_ _03123_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__a21o_1
XANTENNA__05370__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout342_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ _04486_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06516_ _01922_ _02178_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__nor2_1
XANTENNA__07647__B1 _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ _02770_ _03054_ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09235_ net231 _04441_ _04442_ net408 net901 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__a32o_1
X_06447_ _02086_ _02120_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10840__516 vssd1 vssd1 vccd1 vccd1 _10840__516/HI net516 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_118_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04369_ _04384_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__and3_1
X_06378_ _02043_ _02050_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08117_ net761 net760 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05329_ _01008_ _01015_ vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09097_ net212 _04339_ _04340_ net399 net975 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__a32o_1
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07078__A _02726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08048_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[20\]
+ net298 _03577_ vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout88_A _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ clknet_leaf_55_wb_clk_i _00007_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_09999_ clknet_leaf_42_wb_clk_i _00019_ net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07084__Y _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07525__B _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10912_ net657 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_58_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07541__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10843_ net519 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07638__B1 _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10774_ clknet_leaf_65_wb_clk_i _00595_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06157__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05996__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06604__B _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06074__C1 _01760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06613__A1 _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10208_ clknet_leaf_83_wb_clk_i _00212_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_10139_ clknet_leaf_31_wb_clk_i team_07_WB.instance_to_wrap.team_07.recGen.circleDetect
+ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.circlePixel sky130_fd_sc_hd__dfrtp_1
XANTENNA__06129__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05680_ net440 _01376_ vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__xor2_1
XANTENNA__09618__A1 _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06338__Y _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07350_ _02958_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06301_ net438 _01966_ _01968_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06521__A1_N _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07281_ _02915_ _02916_ _00679_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[9\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ _04280_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06232_ _01670_ _01706_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06163_ net114 _01840_ _01843_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__o21a_1
Xhold202 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold213 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05114_ _00826_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
Xhold224 _00466_ vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold235 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\] vssd1 vssd1
+ vccd1 vccd1 net905 sky130_fd_sc_hd__dlygate4sd3_1
X_06094_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[9\] _01776_ vssd1
+ vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__or2_1
Xhold246 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[39\]
+ vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold257 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[5\] vssd1 vssd1
+ vccd1 vccd1 net927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[0\] vssd1 vssd1
+ vccd1 vccd1 net938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _01783_ net153 net740 vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__o21ai_1
X_05045_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[7\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_40_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09853_ _04825_ _04855_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__a21o_1
XANTENNA__06907__A2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout292_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ net195 _04157_ vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__nor2_1
X_09784_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[0\] net269 vssd1
+ vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__or2_1
X_06996_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[11\] _02649_
+ _02651_ _02659_ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__o2bb2a_1
X_08735_ net1166 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ net234 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__mux2_1
XANTENNA__07064__C _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05947_ _01637_ _01640_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout178_X net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _04080_ _04093_ _04084_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07868__B1 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05878_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] _01561_
+ net148 _01571_ _01559_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a32oi_4
X_07617_ _01655_ net169 _03132_ _03172_ _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10324__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08597_ _03623_ _04032_ net139 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07080__B _02209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ _01726_ _03083_ _03085_ _01661_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05894__A2 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07096__A1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07096__B2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07479_ _01618_ _02079_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09218_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10490_ clknet_leaf_15_wb_clk_i _00358_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_09149_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09545__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07571__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ net502 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_45_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05885__A2 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07087__A1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10757_ clknet_leaf_61_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[4\]
+ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07087__B2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10454__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10688_ clknet_leaf_53_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[20\]
+ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06334__B net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07584__B1_N _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06850_ net433 _02520_ _02518_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__a21o_1
XANTENNA__08976__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05801_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] _01486_
+ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__and2_1
XANTENNA__10347__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06781_ _02448_ _02452_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_69_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08520_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[3\] vssd1 vssd1 vccd1 vccd1
+ _03983_ sky130_fd_sc_hd__and3_1
X_05732_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00772_ _00766_
+ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08451_ net469 net475 _03640_ _03657_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05663_ _01374_ _01375_ _01346_ _01366_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[6\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_137_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05413__B _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08382_ net477 _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05594_ _01305_ _01306_ vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07333_ _00675_ _02946_ _02945_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_y\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10195__RESET_B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05700__Y _01413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07264_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__a21o_1
X_09003_ net251 net403 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__mux2_1
X_06215_ net91 _01800_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07195_ _02783_ _02832_ _02845_ _02777_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout305_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06146_ _01823_ _01826_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06077_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__nor2_1
XANTENNA__07356__A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ _01779_ _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05028_ _00753_ _00760_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09836_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__inv_2
XANTENNA__07553__A2 _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ net248 _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__or2_1
X_06979_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\]
+ _02643_ vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08718_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ _04132_ net263 vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__o21ai_1
X_09698_ _04745_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07091__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08649_ _00693_ _04067_ _04059_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_25_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10846__522 vssd1 vssd1 vccd1 vccd1 _10846__522/HI net522 sky130_fd_sc_hd__conb_1
XFILLER_0_37_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10611_ clknet_leaf_49_wb_clk_i _00475_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08266__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10542_ clknet_leaf_20_wb_clk_i _00410_ net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06435__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10473_ clknet_leaf_14_wb_clk_i _00341_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07777__C1 _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06044__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05993__B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11025_ net391 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10933__583 vssd1 vssd1 vccd1 vccd1 _10933__583/HI net583 sky130_fd_sc_hd__conb_1
XANTENNA__07544__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06752__B1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10809_ clknet_leaf_77_wb_clk_i _00630_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_19 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08036__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06283__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06000_ net136 net138 net170 _01687_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__a31o_1
XFILLER_0_113_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05248__X _00961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09509__B1 _04584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ net397 net112 vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06902_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[0\] _02106_ _00749_
+ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a21oi_1
X_07882_ _03329_ _03338_ _03409_ _03436_ _03328_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__o2111a_1
X_11012__640 vssd1 vssd1 vccd1 vccd1 _11012__640/HI net640 sky130_fd_sc_hd__conb_1
XANTENNA__07535__A2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09621_ _04666_ _04690_ _04691_ _04664_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\]
+ vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__a32o_1
X_06833_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\] net174 vssd1 vssd1
+ vccd1 vccd1 _02504_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07904__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07940__C1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ net947 net209 _04655_ vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__o21a_1
X_06764_ net99 _02417_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08503_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[19\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[18\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[20\] _03968_ vssd1 vssd1
+ vccd1 vccd1 _03969_ sky130_fd_sc_hd__nor4_1
X_05715_ net1140 _00797_ _01412_ _01426_ _01427_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__a221o_1
XANTENNA__08496__B1 net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09483_ net977 net206 _04615_ vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__o21a_1
X_06695_ _02284_ _02286_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__nor2_1
XANTENNA__07342__C _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949__590 vssd1 vssd1 vccd1 vccd1 _10949__590/HI net590 sky130_fd_sc_hd__conb_1
XANTENNA_fanout255_A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10376__RESET_B net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ net463 _03561_ _03907_ net477 vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05646_ _01357_ _01358_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_121_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08365_ net461 _03839_ _03840_ _01379_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__o22a_1
X_05577_ _01282_ _01288_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07316_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.nxt_rand_x\[1\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ net460 _03773_ _03675_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07471__A1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07247_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[5\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09566__A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07178_ _01665_ _01724_ _02829_ net205 vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__o211a_2
XFILLER_0_108_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06129_ _01720_ _01735_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_86_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06702__B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout320 net322 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_4
XANTENNA__05785__A1 _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout331 net333 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_4
Xfanout342 net343 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_4
Xfanout353 net357 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_4
Xfanout364 net366 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_4
Xfanout375 net388 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_2
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07814__A _01113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09819_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__and4_1
Xfanout397 _00968_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_4
XANTENNA__07931__C1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07533__B net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05988__B net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput28 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10525_ clknet_leaf_21_wb_clk_i _00393_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput39 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10456_ clknet_leaf_62_wb_clk_i _00016_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07214__A1 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10387_ clknet_leaf_11_wb_clk_i net681 net327 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_23_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05068__X _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05228__B net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11008_ net390 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05244__A team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05500_ net422 _00691_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_16_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06480_ net144 net105 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__nor2_4
XFILLER_0_8_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05431_ _01077_ _01127_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08150_ _03635_ _03636_ vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05362_ net191 _01074_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__or2_1
XANTENNA__06075__A _01748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07101_ _02754_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06506__C _01609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08081_ _00814_ _01429_ net232 net1059 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05293_ net192 _01004_ _01005_ vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__nor3_1
XFILLER_0_71_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07032_ _02251_ _02686_ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06661__C1 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06362__X _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06803__A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07205__A1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07177__Y _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06522__B net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06559__A3 _02232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07934_ _01084_ _03309_ _03316_ net189 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07508__A2 _02262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07865_ _03359_ _03390_ _03288_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09604_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\]
+ _04678_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_3_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06816_ _02484_ _02486_ vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_123_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07796_ net280 _01115_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_123_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[35\]
+ net271 _04647_ net291 net223 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__a221o_1
X_06747_ _02418_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout160_X net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout258_X net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[8\]
+ net272 net293 net221 vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a211o_1
X_06678_ _02184_ _02350_ _02349_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08417_ _00717_ _03891_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__nand2_1
XANTENNA__07692__A1 _03041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05629_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] _01315_
+ _01339_ _01341_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__o211ai_1
X_09397_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[4\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\] vssd1 vssd1
+ vccd1 vccd1 _04555_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ _00126_ _03824_ _03801_ vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06247__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08279_ net469 _03756_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10310_ clknet_leaf_45_wb_clk_i net781 net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_131_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10241_ clknet_leaf_76_wb_clk_i net711 net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_30_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06432__B net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ clknet_leaf_9_wb_clk_i _00182_ net308 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout150 _01567_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_8
Xfanout161 net162 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_4
Xfanout172 _01668_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_4
Xfanout183 _01532_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_4
Xfanout194 _00990_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__buf_2
XANTENNA__06707__B1 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10298__RESET_B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05064__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10227__RESET_B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05999__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07683__A1 _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05446__B1 _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10508_ clknet_leaf_16_wb_clk_i _00376_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06182__X _01863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10439_ clknet_leaf_45_wb_clk_i _00323_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07199__B1 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06342__B net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05980_ net1110 _01633_ _01641_ _01660_ _01673_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[0\]
+ sky130_fd_sc_hd__a2111oi_2
XTAP_TAPCELL_ROW_72_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04931_ net427 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10088__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ net254 _01734_ _02371_ _03114_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06174__B2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06601_ net123 _01652_ _02014_ net158 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a211o_1
XANTENNA__07910__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ net131 net138 _01719_ _01903_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__a31o_1
X_09320_ _00661_ _04500_ net228 vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06532_ _02188_ _02199_ _02205_ _02183_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__or4b_1
XANTENNA__06357__X _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09251_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ _04449_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07674__A1 _02055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06463_ _02053_ _02136_ _02135_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06517__B _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08202_ net462 _01383_ _03680_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05414_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] _01062_ vssd1
+ vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__nand2_1
X_09182_ net211 _04401_ _04402_ net400 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_32_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06394_ _01693_ _01696_ _02052_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08133_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[17\]
+ _03619_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05345_ net437 _01048_ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout120_A _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout218_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ net396 net298 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ _03585_ vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__a221o_1
XFILLER_0_102_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05276_ net427 _00983_ _00670_ vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07015_ _02671_ vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08966_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[6\] net813
+ net447 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07917_ net277 _03354_ _03363_ net275 vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__o22a_1
X_08897_ _00708_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[5\]
+ net481 vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07848_ _01679_ _03380_ _03388_ _01689_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07901__A2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07779_ net435 net112 _03275_ _03333_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09518_ net896 net207 _04636_ vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__o21a_1
XANTENNA__07811__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10790_ clknet_leaf_77_wb_clk_i _00611_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07665__A1 _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09449_ _01415_ _04589_ _04586_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06427__B net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08614__B1 _00960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07968__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05979__A1 _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10224_ clknet_leaf_85_wb_clk_i _00228_ net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10155_ clknet_leaf_2_wb_clk_i team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10086_ clknet_leaf_69_wb_clk_i _00144_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[10\]
+ vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10988_ net629 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_128_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05522__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06337__B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05130_ _00835_ _00841_ _00842_ vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07959__A2 _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08044__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold406 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[1\] vssd1 vssd1 vccd1
+ vccd1 net1076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold417 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[1\] vssd1
+ vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold428 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\] vssd1 vssd1 vccd1
+ vccd1 net1098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold439 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\] vssd1 vssd1
+ vccd1 vccd1 net1109 sky130_fd_sc_hd__dlygate4sd3_1
X_05061_ _00790_ vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_74_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09030__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[13\] _01448_
+ _04160_ net864 vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__o31ai_1
X_08751_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[25\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ net234 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__mux2_1
X_05963_ net218 net199 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__nor2_4
XFILLER_0_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04914_ net938 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
X_07702_ net86 _01635_ _03257_ _03255_ _03251_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__o311a_1
XFILLER_0_75_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08682_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ _04082_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__nor2_1
X_05894_ _01574_ _01575_ _00715_ _01569_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_36_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07633_ _01660_ _02167_ _03080_ _03117_ _03190_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__a41o_1
XFILLER_0_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout168_A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07190__Y _02842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07564_ net102 _03078_ _03121_ _03122_ _01646_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__a2111o_1
X_09303_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ _04486_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__a21o_1
X_06515_ _02054_ _02115_ _02155_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07647__A1 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07495_ _00685_ _00941_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout335_A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09234_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04435_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05151__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06446_ net168 _02069_ _02088_ _02110_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09165_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04384_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06377_ _02050_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout123_X net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08116_ net747 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[6\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05328_ _01008_ _01015_ vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09096_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ _04337_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08047_ net452 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[18\]
+ net394 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06622__A2 _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05259_ _00671_ net429 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04989__Y _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09572__A1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06386__A1 _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07806__B net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ clknet_leaf_45_wb_clk_i _00001_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07583__B1 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ net491 _04241_ vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__and2b_1
XANTENNA__07822__A _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10911_ net656 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XFILLER_0_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07541__B _02048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ net518 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__06438__A _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05342__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08835__B1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ clknet_leaf_65_wb_clk_i _00594_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05996__B net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06074__B1 _01759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10207_ clknet_leaf_81_wb_clk_i _00211_ net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10138_ clknet_leaf_31_wb_clk_i team_07_WB.instance_to_wrap.team_07.borderGen.synchronized_rectangle_pixel
+ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.borderGen.borderPixel
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06129__A1 _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10069_ clknet_leaf_35_wb_clk_i _00127_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09866__A2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07451__B net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08039__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05252__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10863__539 vssd1 vssd1 vccd1 vccd1 _10863__539/HI net539 sky130_fd_sc_hd__conb_1
XFILLER_0_45_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06300_ net187 _01975_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_98_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07280_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[9\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06231_ _01892_ _01895_ _01896_ _01909_ _01889_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a41o_1
XFILLER_0_116_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06852__A2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06162_ net120 _01797_ _01804_ _01840_ net114 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__a32o_1
Xhold203 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[3\] vssd1 vssd1
+ vccd1 vccd1 net873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold214 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__dlygate4sd3_1
X_05113_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[1\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[2\] vssd1 vssd1 vccd1
+ vccd1 _00826_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_113_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold225 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[15\]
+ vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__dlygate4sd3_1
X_06093_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[7\]
+ _01775_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__or3_1
Xhold236 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[26\]
+ vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold247 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[0\]
+ vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[10\]
+ vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _01783_ _04870_ _04900_ vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__o21ai_1
X_05044_ _00652_ _00775_ _00763_ vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__o21ai_1
Xhold269 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[29\]
+ vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07907__A _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09852_ net269 _04854_ _04856_ net247 net1038 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__a32o_1
X_08803_ net1168 _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__xor2_1
X_09783_ net269 _04807_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nand2b_2
X_06995_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[12\] _02650_
+ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout285_A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ net1162 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[8\]
+ net238 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__mux2_1
X_05946_ net98 net88 net276 _01638_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__a31o_1
XANTENNA__07868__A1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04047_ _04072_ _04089_ _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__o311a_1
X_05877_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _01555_
+ _01546_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout452_A team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__B _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07616_ net126 _01676_ _03173_ _02262_ net167 vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__a32o_1
X_08596_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[20\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\] _03621_
+ net863 vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__o31ai_1
XANTENNA__06258__A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout240_X net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07547_ _03105_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07096__A2 _01921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07478_ _01626_ _01635_ _02176_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__or3b_1
XANTENNA__08293__A1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ net230 _04428_ _04429_ net406 net996 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_20_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06429_ _01722_ _02056_ _02054_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07089__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ net210 _04377_ _04378_ net399 net991 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__a32o_1
XANTENNA__09242__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10769__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06056__B1 _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09079_ net213 _04326_ _04327_ net400 net999 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07817__A _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05583__C_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07308__B1 _02930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ net501 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_45_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10299__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ clknet_leaf_66_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[3\]
+ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06455__X _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10687_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[19\]
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_93_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06631__A _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05800_ _01490_ _01493_ _01491_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__and4bb_1
X_06780_ _00984_ net174 _02451_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_69_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05731_ _00709_ _00710_ _01436_ _01434_ net486 vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a32o_1
XFILLER_0_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08450_ _03662_ _03815_ _03922_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__o211a_1
X_05662_ _01255_ _01257_ _01278_ _01323_ _00679_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_106_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07401_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\] _02992_
+ net480 vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08381_ _03856_ team_07_WB.instance_to_wrap.team_07.defusedGen.defusedPixel team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__mux2_2
XFILLER_0_133_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05593_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] vssd1 vssd1 vccd1
+ vccd1 _01306_ sky130_fd_sc_hd__or3b_2
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07332_ net431 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09472__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07263_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06214_ _01807_ _01892_ _01893_ _01820_ _01891_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a221o_1
X_09002_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ net2 _04252_ _04269_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__a211oi_1
X_07194_ _02845_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06145_ net91 _01803_ _01825_ net101 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_41_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout200_A _01517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06076_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[6\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\] vssd1 vssd1 vccd1
+ vccd1 _01763_ sky130_fd_sc_hd__and3b_1
XANTENNA__10164__RESET_B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09904_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[12\] _01778_
+ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05027_ net287 _00751_ vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input5_A gpio_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ _04840_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout190_X net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09766_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\] _04790_ _04767_
+ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a21boi_1
X_06978_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _02643_
+ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__xor2_1
X_08717_ _04128_ _04130_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__nor2_1
X_05929_ net284 net275 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09697_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\]
+ net250 _04742_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06259__Y _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08648_ _04054_ _04075_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__a21o_1
XANTENNA__06513__A1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10885__561 vssd1 vssd1 vccd1 vccd1 _10885__561/HI net561 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_25_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[16\]
+ _03618_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__nand2_1
X_10610_ clknet_leaf_49_wb_clk_i net924 net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ clknet_leaf_20_wb_clk_i _00409_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10472_ clknet_leaf_14_wb_clk_i _00340_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06029__B1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07777__B1 _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07529__B1 _02110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05067__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ net644 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XANTENNA__05354__X _01067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07701__B1 _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10808_ clknet_leaf_77_wb_clk_i _00629_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10739_ clknet_leaf_72_wb_clk_i _00569_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10675__RESET_B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09937__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07950_ _03471_ _03472_ _03503_ _03504_ _03502_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06901_ _02527_ _02542_ _02570_ _02571_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a22o_1
X_07881_ _03417_ _03418_ _03434_ _03435_ _03412_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09620_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[14\] _04688_ vssd1
+ vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__nand2_1
XANTENNA__07535__A3 _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06832_ _02501_ _02502_ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_108_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912__657 vssd1 vssd1 vccd1 vccd1 net657 _10912__657/LO sky130_fd_sc_hd__conb_1
X_09551_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[44\]
+ net273 net293 net225 vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a211o_1
X_10869__545 vssd1 vssd1 vccd1 vccd1 _10869__545/HI net545 sky130_fd_sc_hd__conb_1
X_06763_ _02425_ _02431_ _02434_ _02423_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_125_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08502_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[17\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[16\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__or4b_1
X_05714_ net414 _00827_ _01423_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__nor3_1
XFILLER_0_77_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08496__A1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06694_ _01624_ net84 _02313_ net253 _02366_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a221o_1
X_09482_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[15\]
+ net270 _04612_ _04614_ net223 vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08433_ net465 _03857_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05645_ net419 _00676_ _00677_ _01356_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_121_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08364_ _03678_ _03731_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__or2_1
X_05576_ _01282_ _01288_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__nand2_1
XANTENNA__06536__A _02178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05440__A _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07315_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[1\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08295_ net419 _03678_ _03772_ net461 vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout415_A _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07246_ _00720_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ _02894_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[3\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07177_ net205 _02828_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__nand2_2
XFILLER_0_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout203_X net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06128_ net289 net107 net105 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__or3_1
XANTENNA__06271__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06702__C _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06059_ net946 _01633_ _01746_ _01747_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[5\]
+ sky130_fd_sc_hd__a211oi_2
Xfanout310 net312 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_4
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout332 net333 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout343 net389 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_4
Xfanout354 net357 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_2
Xfanout365 net366 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_4
Xfanout376 net378 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_4
Xfanout387 net388 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_2
X_09818_ net1135 _04830_ _04831_ _04832_ vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__o22a_1
Xfanout398 _00943_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_2
XANTENNA__07814__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09749_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\] _04777_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__a21o_1
XANTENNA__07533__C net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08487__A1 _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08645__B _04070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
X_10524_ clknet_leaf_20_wb_clk_i _00392_ net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10086__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput29 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06670__B1 _02027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10455_ clknet_leaf_62_wb_clk_i _00015_ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_122_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08411__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10386_ clknet_leaf_11_wb_clk_i net682 net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_62_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ net390 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06725__B2 _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output44_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10981__622 vssd1 vssd1 vccd1 vccd1 _10981__622/HI net622 sky130_fd_sc_hd__conb_1
XANTENNA__07740__A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05430_ _01026_ _01110_ _01106_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06356__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05361_ _01005_ _01019_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06075__B _01761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07100_ _02726_ _02729_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__and2b_1
X_08080_ _03591_ _03592_ _00815_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__mux2_1
XANTENNA__07453__A2 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05292_ _00675_ _00998_ vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__nand2_2
XFILLER_0_114_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07031_ net265 net83 _02335_ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06803__B team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06522__C _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06413__B1 _02086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08982_ _00664_ _04249_ _04250_ _04251_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__a31oi_1
X_07933_ _03305_ _03442_ _03444_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07864_ _03352_ _03360_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__nand2b_1
XANTENNA__06716__A1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[8\] _04678_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a21o_1
X_06815_ net286 net434 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_123_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07795_ _03348_ _03349_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_123_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05154__B _00863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ _00666_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\] vssd1 vssd1
+ vccd1 vccd1 _04647_ sky130_fd_sc_hd__a21oi_1
X_06746_ _00670_ _00983_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__xnor2_2
X_09465_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[8\]
+ net221 _04605_ net909 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__a22o_1
X_06677_ _01636_ net84 _02250_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__a21oi_1
X_08416_ net469 net471 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__and2b_1
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05628_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] net443
+ team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\] _01338_ _01340_ vssd1
+ vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__o311a_1
XFILLER_0_65_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09396_ net414 net417 _01475_ _04554_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__o31a_1
XFILLER_0_114_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08347_ _03753_ _03814_ _03818_ _03823_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05559_ _01269_ _01271_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08278_ _03638_ _03641_ _03755_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__or3_1
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07229_ _02860_ _02856_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10240_ clknet_leaf_82_wb_clk_i net687 net321 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10171_ clknet_leaf_10_wb_clk_i _00181_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout140 _03625_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
Xfanout151 _04869_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_2
Xfanout162 net163 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_4
Xfanout173 _01543_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_8
XANTENNA__06707__A1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout184 net186 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_8
Xfanout195 net196 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_2
XANTENNA__05345__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10965__606 vssd1 vssd1 vccd1 vccd1 _10965__606/HI net606 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_83_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05064__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07560__A _03117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05999__B net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05351__Y _01064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07683__A2 _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05080__A team_07_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10507_ clknet_leaf_16_wb_clk_i _00375_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07772__A1_N _01688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05667__C_N team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10438_ clknet_leaf_45_wb_clk_i _00322_ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07199__A1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10369_ clknet_leaf_23_wb_clk_i net691 net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06061__D _00961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_04930_ net426 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
XANTENNA__05255__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06174__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06600_ _01804_ _02013_ net254 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__a21o_1
X_07580_ _03136_ _03138_ _03129_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05921__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06531_ _01624_ _02166_ net84 _02204_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_0_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09250_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[10\]
+ _04449_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__a21o_1
X_06462_ net104 net166 _02104_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07674__A2 _02282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08201_ net420 net462 _01257_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__and3b_1
XFILLER_0_84_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05413_ _01047_ _01109_ _01121_ _01125_ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__and4b_1
X_09181_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ _04399_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06393_ _00649_ _02065_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_32_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08132_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[16\]
+ _03618_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__or2_1
X_05344_ _00668_ _01056_ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__nor2_4
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06634__B1 _02178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ net456 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__and2b_1
XFILLER_0_109_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05275_ _00979_ _00987_ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__nand2_2
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout113_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07014_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.idle team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.internalSck
+ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__and2b_2
XFILLER_0_114_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10918__663 vssd1 vssd1 vccd1 vccd1 net663 _10918__663/LO sky130_fd_sc_hd__conb_1
X_08965_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[5\] net842
+ net447 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout482_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ _03455_ _03461_ _03466_ _03470_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__a22oi_1
X_08896_ _04213_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[5\]
+ _04209_ vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__mux2_1
XANTENNA__09887__B1 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07847_ net274 _03392_ _03401_ _03398_ _03393_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__o32a_1
X_07778_ net435 net112 _03330_ _03332_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09517_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[29\]
+ net271 net292 _04582_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06729_ _02079_ _02149_ _02375_ _02066_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09448_ net930 net208 _04594_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__o21a_1
XANTENNA__05612__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07665__A2 _02055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08862__A1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09379_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ _04541_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06724__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05979__A2 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10223_ clknet_leaf_86_wb_clk_i _00227_ net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06928__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input43_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10154_ clknet_leaf_1_wb_clk_i net846 net308 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[5\]
+ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ clknet_leaf_69_wb_clk_i _00143_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10987_ net628 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05081__Y team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08853__A1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07959__A3 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold407 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold418 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[4\] vssd1 vssd1
+ vccd1 vccd1 net1088 sky130_fd_sc_hd__dlygate4sd3_1
X_05060_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\] _00788_ vssd1
+ vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09945__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold429 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[17\] vssd1 vssd1
+ vccd1 vccd1 net1099 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07041__B1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08750_ net1150 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__mux2_1
X_05962_ net199 _01645_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__nand2_1
X_07701_ net111 _01921_ _02176_ _02332_ _02216_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__a221o_1
X_04913_ net851 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
X_08681_ _04034_ _04083_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05893_ _01586_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07632_ _01632_ _02182_ _03189_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__and3b_1
XFILLER_0_36_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05713__A _01413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07563_ _01543_ _01701_ _02743_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__and3_1
X_09302_ net229 _04488_ _04489_ net404 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06514_ _01711_ _02047_ _02184_ _02187_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__a31o_1
XANTENNA__07647__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07494_ net283 _00749_ net119 net89 vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__a31o_1
X_09233_ _04440_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06445_ net281 net284 net268 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_118_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout328_A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09164_ net1122 net401 net210 _04389_ vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06376_ _02047_ _02049_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__and2_2
XFILLER_0_72_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08115_ net765 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05327_ _01039_ vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
X_09095_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[6\]
+ _04337_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout116_X net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ _03576_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[17\]
+ net456 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__mux2_1
X_05258_ net428 _00672_ vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05189_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00901_ vssd1 vssd1
+ vccd1 vccd1 _00902_ sky130_fd_sc_hd__or2_1
X_09997_ clknet_leaf_41_wb_clk_i _00018_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06386__A2 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__A1 _01655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08948_ _00709_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_col _04234_
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_cleared vssd1 vssd1 vccd1 vccd1
+ _04241_ sky130_fd_sc_hd__a31o_1
X_08879_ _01109_ _04198_ _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__a21oi_1
X_10910_ net655 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XANTENNA__07822__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ net517 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_67_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06438__B _02110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10772_ clknet_leaf_66_wb_clk_i _00593_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07638__A2 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06454__A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06460__Y _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10206_ clknet_leaf_83_wb_clk_i _00210_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07574__A1 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07574__B2 _02836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ clknet_leaf_31_wb_clk_i team_07_WB.instance_to_wrap.team_07.recMOD.modHighlightDetect
+ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.modHighlightPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10068_ clknet_leaf_35_wb_clk_i _00126_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ sky130_fd_sc_hd__dfxtp_4
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06129__A2 _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06629__A _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05252__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06230_ _01821_ _01890_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06161_ net114 _01840_ _01841_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07894__S net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05112_ net990 _00817_ _00823_ net1018 vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__a22o_1
Xhold204 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06092_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[6\] _01774_ vssd1
+ vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__or2_1
Xhold215 team_07_WB.instance_to_wrap.team_07.label_num_bus\[0\] vssd1 vssd1 vccd1
+ vccd1 net885 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold226 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[30\]
+ vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold237 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[42\]
+ vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09920_ _01782_ net153 net738 vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__o21ai_1
X_05043_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\]
+ _00773_ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__and3_1
Xhold248 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[28\]
+ vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold259 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[19\]
+ vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07907__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09554__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09851_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08802_ _04155_ _04156_ net195 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__a21oi_1
X_09782_ _00655_ _00656_ _00764_ _04806_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a41o_1
X_06994_ _02652_ _02657_ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06773__C1 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ net1073 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ net234 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__mux2_1
X_05945_ net98 net89 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__nand2_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout278_A _00651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ _04085_ _04090_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__a22oi_2
X_05876_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] _01561_
+ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__nand2_1
XANTENNA__07868__A2 _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06539__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07615_ _02873_ _03120_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__nand2_1
XANTENNA__08457__C _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08595_ _03622_ _04031_ net146 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__o21a_1
XANTENNA__06258__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07546_ _02235_ _02734_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07477_ net266 _01619_ _02779_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09216_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06428_ _01722_ _02056_ _02054_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_20_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06274__A _00684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09147_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__or2_1
X_06359_ _01689_ _01936_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__nor2_2
XANTENNA__07089__B _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06056__A1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08029_ net413 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ net294 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ _03565_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__a221o_1
XANTENNA__07817__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout93_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09545__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__A1 _02235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10824_ net500 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_45_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10755_ clknet_leaf_66_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[2\]
+ net352 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10686_ clknet_leaf_52_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[18\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06184__A net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06912__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06350__C net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10830__506 vssd1 vssd1 vccd1 vccd1 _10830__506/HI net506 sky130_fd_sc_hd__conb_1
XFILLER_0_101_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05730_ _00711_ _01435_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06359__A _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05661_ _01300_ _01373_ _01278_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07400_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[5\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[6\]
+ _02990_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08380_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.boomGen.boomPixel vssd1 vssd1 vccd1 vccd1 _03856_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_92_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05592_ net421 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\] vssd1 vssd1 vccd1
+ vccd1 _01305_ sky130_fd_sc_hd__or3b_2
XFILLER_0_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07331_ _00965_ _01175_ _01190_ _01192_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07262_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09001_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ net2 net334 vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06213_ _01805_ _01807_ _01890_ _01892_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__and4bb_1
XANTENNA__09676__Y _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07193_ _02822_ _02826_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06144_ _01802_ _01824_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__xor2_1
XANTENNA__06822__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06075_ _01748_ _01761_ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09903_ net850 net154 net151 _04889_ vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__a22o_1
X_05026_ net266 _00759_ vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout395_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05157__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09834_ net269 _04842_ _04843_ net247 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__a32o_1
X_09765_ _04767_ _04791_ _04792_ net249 net1055 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__a32o_1
XFILLER_0_77_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06977_ _02643_ _02644_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout183_X net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06761__A2 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ _04131_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ _04128_ vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__mux2_1
X_05928_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] net288
+ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__or2_1
X_09696_ _00700_ _04730_ _04743_ _04744_ _04734_ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__o311a_1
XFILLER_0_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08647_ _04058_ _04060_ _04074_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__and3b_1
XFILLER_0_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05859_ _01548_ _01550_ _01551_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06513__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ _03997_ _04022_ _03996_ vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07529_ net170 net104 _02110_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08266__A2 _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ clknet_leaf_21_wb_clk_i _00408_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10471_ clknet_leaf_14_wb_clk_i _00339_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06029__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07777__B2 _01104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout96_X net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11023_ net391 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05067__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__A _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05960__B1 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07162__C1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07701__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07701__B2 _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05370__X _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ clknet_leaf_77_wb_clk_i _00628_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07465__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10738_ clknet_leaf_60_wb_clk_i _00568_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10669_ clknet_leaf_64_wb_clk_i net952 net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08841__B _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07217__B1 _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06440__A1 _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06900_ net268 _02568_ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__or2_1
X_07880_ net106 _03381_ _03387_ _01692_ _03380_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__o32a_1
X_06831_ net160 _02500_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_108_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07940__A1 _01067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ net960 net209 _04654_ vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__o21a_1
X_06762_ _02424_ _02425_ _02433_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__nor3_1
X_08501_ team_07_WB.instance_to_wrap.team_07.audio_0.bm_state\[1\] _00657_ vssd1 vssd1
+ vccd1 vccd1 _03967_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_125_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05713_ _01413_ _01424_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09481_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ _04613_ net291 vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__o21a_1
X_06693_ _02209_ _02259_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08432_ _03631_ _03637_ _03901_ _03905_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_19_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05644_ net419 _01356_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\] vssd1 vssd1 vccd1
+ vccd1 _01357_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_37_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08363_ _01256_ _03729_ _03838_ net462 vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__o22a_1
X_05575_ _01286_ _01287_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06536__B _02209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07314_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ net770 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ _00722_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_y\[2\]
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_116_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08294_ net462 _03771_ _03680_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07245_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout310_A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout408_A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07208__B1 _00943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07176_ net187 _01901_ net199 vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07759__A1 _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06127_ net287 _01720_ _01735_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06058_ _01641_ _01738_ _01744_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__or3_1
Xfanout300 _00942_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout311 net312 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_4
Xfanout322 net323 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05009_ net42 net40 net43 _00744_ vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__and4_1
Xfanout333 net338 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_2
Xfanout344 net346 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_4
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_4
Xfanout366 net375 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_4
X_09817_ _00657_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[3\] vssd1
+ vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__nor2_1
Xfanout377 net378 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_4
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__clkbuf_4
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_2
XFILLER_0_119_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09748_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[7\]
+ _04777_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__nand3_1
XFILLER_0_119_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09679_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _04704_ vssd1
+ vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08645__C _04071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_66_wb_clk_i_X clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08942__A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10523_ clknet_leaf_20_wb_clk_i _00391_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput19 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06670__A1 _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ clknet_leaf_31_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing_mod_locator.nxt_mod_row
+ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10385_ clknet_leaf_11_wb_clk_i net705 net326 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_20_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06973__A2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11006_ net390 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06186__B1 _01863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07686__B1 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05697__C1 _00962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06356__B net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05360_ net194 _01004_ _01010_ _01071_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__or4_1
XFILLER_0_82_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05291_ _00993_ _00995_ vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__or2_4
XFILLER_0_70_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07030_ net129 _01677_ _01708_ _02684_ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__or4_1
XANTENNA__06661__A1 _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06372__A _01642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06661__B2 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06413__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10836__512 vssd1 vssd1 vccd1 vccd1 _10836__512/HI net512 sky130_fd_sc_hd__conb_1
X_08981_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__nand3_1
X_07932_ _03311_ _03324_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_127_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07863_ _01650_ _03321_ _03326_ _01692_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06716__A2 _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__A1 _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09602_ net1094 _04678_ vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__xor2_1
X_06814_ net280 net434 _02484_ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07794_ net282 _01069_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_123_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09533_ net937 net206 _04646_ vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06745_ _00673_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ _02409_ _02416_ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout260_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07677__B1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[7\]
+ net221 _04605_ net893 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06676_ _01639_ _02348_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__and2_1
XANTENNA__06547__A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08415_ _03646_ _03889_ _03657_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__a21oi_1
X_05627_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] _01319_
+ _01328_ net421 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__o22a_1
X_09395_ _01425_ _04551_ _04553_ net233 vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08346_ _03657_ _03820_ _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__o21ai_1
X_05558_ _01254_ _01268_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08277_ net470 _00717_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__nor2_1
X_05489_ _00688_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07228_ _02081_ _02775_ _02877_ _02878_ _02767_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__a32o_1
XFILLER_0_61_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06652__A1 _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06282__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08929__A0 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07159_ _02065_ net81 _02736_ _02807_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__a22o_1
X_10893__650 vssd1 vssd1 vccd1 vccd1 net650 _10893__650/LO sky130_fd_sc_hd__conb_1
XFILLER_0_121_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10170_ clknet_leaf_10_wb_clk_i _00180_ net324 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout130 _03653_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
XFILLER_0_100_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout141 net143 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_4
Xfanout152 _04869_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout163 _01557_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__buf_4
Xfanout174 net180 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_4
Xfanout185 net186 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06707__A2 _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 _04144_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_83_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08937__A _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07668__B1 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07560__B _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05361__A _01005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06340__B1 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07683__A3 _01935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08093__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07559__Y _03118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06643__A1 _02031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10506_ clknet_leaf_14_wb_clk_i _00374_ net332 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10236__RESET_B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06192__A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10437_ clknet_leaf_44_wb_clk_i _00321_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07199__A2 _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ clknet_leaf_22_wb_clk_i net722 net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06920__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__B _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10299_ clknet_leaf_54_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[12\]
+ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05255__B team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05823__X _01517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06530_ _02202_ _02203_ _01618_ _02164_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06367__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07123__A2 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08320__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06461_ net267 _00755_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__or2_2
X_08200_ net419 _03678_ _03677_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05412_ _01054_ _01117_ _01122_ _01124_ vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__and4b_1
X_09180_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[11\]
+ _04399_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06392_ net286 net283 _01621_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__and3_2
XFILLER_0_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06654__X _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08131_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[15\]
+ _03617_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05343_ net437 _00669_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__nand2_4
XANTENNA__06373__Y _02047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08062_ net981 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ net296 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__mux2_1
X_05274_ net426 _00984_ _00983_ vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07013_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.idle
+ vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_116_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout106_A _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__A1 _03753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06830__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08964_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] net829
+ net447 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__mux2_1
X_07915_ net256 _03376_ _03469_ _03468_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__a31o_1
X_08895_ _00708_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[4\]
+ net481 vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__o21a_1
X_10988__629 vssd1 vssd1 vccd1 vccd1 _10988__629/HI net629 sky130_fd_sc_hd__conb_1
XANTENNA__05165__B _00860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ _03345_ _03395_ _03399_ _03400_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__nand4_1
XFILLER_0_98_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07661__A _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ _00669_ net118 _02212_ _01104_ _02191_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__a221o_1
XANTENNA__06570__B1 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04989_ net466 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
X_06728_ net265 _02149_ _02375_ _02134_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a22oi_1
X_09516_ net939 net207 _04635_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09447_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[1\]
+ net272 _04593_ net290 net220 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06659_ net279 _02331_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__or2_4
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08862__A2 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09378_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ _04541_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08329_ net461 _03727_ _03728_ _03732_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__o31a_1
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10222_ clknet_leaf_84_wb_clk_i _00226_ net316 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10153_ clknet_leaf_2_wb_clk_i net734 net308 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07050__B2 _02699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10084_ clknet_leaf_69_wb_clk_i _00142_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input36_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[7\]
+ vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10986_ net627 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_58_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10488__RESET_B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08853__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06474__X _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06915__A _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07813__B1 _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold408 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[10\] vssd1 vssd1
+ vccd1 vccd1 net1078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.tft_reset vssd1 vssd1 vccd1
+ vccd1 net1089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07041__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05961_ net126 _01654_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__nor2_4
X_07700_ net265 _01627_ _02150_ _03250_ _03252_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__o311a_1
X_04912_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _00652_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08680_ _04103_ _04104_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__a21o_1
X_05892_ _01561_ _01568_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__xor2_2
X_07631_ _01708_ _02263_ _03188_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07481__A _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07562_ _01740_ _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09301_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ _04486_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06513_ net87 net84 _02186_ _01660_ _02079_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07493_ _02128_ net83 _03052_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09232_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04435_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__and3_1
X_06444_ _02084_ _02114_ _02117_ _02109_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__o31a_1
XFILLER_0_91_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09163_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[6\]
+ _04388_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_118_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06375_ net188 net181 _02048_ _01684_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout223_A _04582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08114_ net773 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[4\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05326_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_x\[0\]
+ _00984_ _00985_ vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__o21a_1
X_09094_ net212 _04336_ _04338_ net399 net1116 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08045_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[19\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ net452 vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__mux2_1
X_05257_ net435 net397 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__nand2_2
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07656__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05188_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[25\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[27\]
+ team_07_WB.instance_to_wrap.team_07.label_num_bus\[29\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[31\]
+ _00899_ _00900_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__mux4_2
X_09996_ clknet_leaf_40_wb_clk_i _00035_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09871__A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ net490 _04240_ vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__and2b_1
XANTENNA__10232__D net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08878_ _04199_ _04200_ _04202_ _00964_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__o31a_1
X_07829_ _01058_ net216 net197 _01095_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__a22o_1
X_10840_ net516 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_6_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05897__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10771_ clknet_leaf_66_wb_clk_i _00592_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07023__A1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ clknet_leaf_86_wb_clk_i _00209_ net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07023__B2 team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07574__A2 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10136_ clknet_leaf_31_wb_clk_i team_07_WB.instance_to_wrap.team_07.recMOD.modSquaresDetect
+ net359 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.modSquaresPixel
+ sky130_fd_sc_hd__dfrtp_1
X_10067_ clknet_leaf_28_wb_clk_i _00125_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.frameBufferLowNibble
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10642__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload1_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10969_ net610 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10251__RESET_B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06364__B _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06160_ net114 _01840_ _01807_ _01805_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08860__A _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05111_ net1049 _00824_ _00825_ net1018 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__a22o_1
Xhold205 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[20\] vssd1 vssd1
+ vccd1 vccd1 net875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06091_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[4\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[5\]
+ _01773_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_113_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold216 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[23\]
+ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _00490_ vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\] vssd1 vssd1
+ vccd1 vccd1 net908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05042_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[4\] _00773_ vssd1
+ vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__nand2_1
Xhold249 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[3\]
+ vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold44_A team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08071__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[13\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[12\]
+ _04850_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08801_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[7\] _04154_ vssd1
+ vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__or2_1
X_06993_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[13\] _02651_
+ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__or2_1
X_09781_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\] _00654_ vssd1
+ vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06773__B1 _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08732_ net1051 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__mux2_1
X_05944_ net95 net93 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__nor2_1
XANTENNA__09711__B1 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ _04049_ _04050_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ _04086_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__o221a_1
X_05875_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] net147
+ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__xnor2_4
XANTENNA__06539__B _02212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07868__A3 _02106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout173_A _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07614_ net104 net164 _03134_ _03171_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__a211o_1
XANTENNA__05879__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08594_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\]
+ _03621_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07545_ _03098_ _03099_ _03103_ net166 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout340_A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07476_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.internalSck team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.cs
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sck
+ sky130_fd_sc_hd__and2_1
XFILLER_0_9_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09215_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06427_ net280 net283 _00045_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09146_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06358_ _02031_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06056__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05309_ _01021_ vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09077_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06289_ net441 net132 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06561__Y _02235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08028_ net453 net451 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_49_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout86_A _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ clknet_leaf_83_wb_clk_i _00084_ net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07325__S _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06531__A3 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10823_ net499 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_138_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06819__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10754_ clknet_leaf_66_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[1\]
+ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06465__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10685_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[17\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06184__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06350__D _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10119_ clknet_leaf_27_wb_clk_i _00157_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06359__B _01936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05660_ _01369_ _01372_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__nor2_1
XANTENNA__05263__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10432__RESET_B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05591_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[14\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] vssd1 vssd1 vccd1
+ vccd1 _01304_ sky130_fd_sc_hd__or3b_2
XFILLER_0_58_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07330_ _02942_ _02944_ _02936_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.next_pos_x\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09472__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07483__A1 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07261_ _00718_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[9\]
+ _02903_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[9\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08680__B1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09000_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ net1 _04268_ vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06212_ net110 _01801_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07192_ _02830_ _02833_ _02843_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06143_ net218 _01799_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06381__Y _02055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06074_ _01395_ _01408_ _01759_ _01760_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__o211a_1
X_09902_ _01778_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05025_ net284 _00753_ vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__or2_4
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09833_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\] _04840_ vssd1
+ vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout290_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09764_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\]
+ _04783_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\] vssd1 vssd1
+ vccd1 vccd1 _04792_ sky130_fd_sc_hd__a31o_1
X_06976_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] _02641_
+ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08715_ net263 _01756_ _04130_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__and3_1
X_05927_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] net288
+ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__nor2_2
X_09695_ net250 _04742_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout176_X net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08646_ _01475_ _01480_ _04070_ net478 vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__o211a_4
XFILLER_0_95_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05858_ _01550_ _01551_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07710__A2 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10102__RESET_B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08577_ _03618_ _04021_ net139 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05789_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row net418 _01436_
+ _01434_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\] vssd1
+ vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__a32o_1
XANTENNA__06556__Y _02230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ net102 _03079_ _03082_ net156 vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07459_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ net395 net296 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ _03030_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[7\]
+ sky130_fd_sc_hd__a221o_1
XANTENNA__08671__B1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10470_ clknet_leaf_20_wb_clk_i _00338_ net337 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.debounce
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06029__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09129_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ net332 _04358_ net1130 vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__a41o_1
XFILLER_0_115_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05237__B1 team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07777__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05788__A1 _00709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05348__B _01000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10853__529 vssd1 vssd1 vccd1 vccd1 _10853__529/HI net529 sky130_fd_sc_hd__conb_1
XANTENNA__07529__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11022_ net391 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout89_X net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05916__X _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07934__C1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05364__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05960__A1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07162__B1 _02767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07701__A2 _01921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ clknet_leaf_78_wb_clk_i _00627_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07465__A1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10737_ clknet_leaf_79_wb_clk_i _00567_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_132_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10668_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[0\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07217__A1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10599_ clknet_leaf_54_wb_clk_i _00463_ net367 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06830_ net160 _02500_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_108_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07940__A2 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06761_ _00973_ net201 _02430_ _02432_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08500_ _00656_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] vssd1
+ vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__nor2_1
X_05712_ _01424_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06692_ net175 _01722_ _02014_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__a21oi_2
X_09480_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\] vssd1
+ vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_78_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08431_ _03663_ _03903_ _03904_ _00703_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05643_ _01354_ _01355_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08362_ _00730_ _01258_ _03725_ _03837_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__o31a_1
XFILLER_0_92_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05574_ _01284_ _01285_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07313_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ net1186 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.nxt_rand_x\[1\]
+ sky130_fd_sc_hd__and2b_1
X_08293_ net421 _00730_ _01258_ _03687_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__o31a_1
XFILLER_0_18_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07244_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07175_ _02822_ _02826_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06126_ _01797_ _01804_ net117 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09976__SET_B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06057_ _01644_ _01739_ _01741_ _01745_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__a31o_1
X_10956__597 vssd1 vssd1 vccd1 vccd1 _10956__597/HI net597 sky130_fd_sc_hd__conb_1
Xfanout301 _00831_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_4
X_05008_ net75 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
Xfanout312 net323 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_2
Xfanout323 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_2
Xfanout334 net335 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 net346 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_4
Xfanout356 net357 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_4
X_09816_ _04829_ _04831_ vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__and2_1
Xfanout367 net375 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_4
Xfanout378 net381 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__buf_2
Xfanout389 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10354__RESET_B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07392__B1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ _04779_ _04778_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06959_ _02608_ _02611_ _02629_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08495__A _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\] _04729_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07695__A1 _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[4\]
+ _04051_ _04056_ _00707_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_64_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10522_ clknet_leaf_20_wb_clk_i _00390_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10453_ clknet_leaf_57_wb_clk_i team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing_mod_locator.nxt_mod_col
+ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_col
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10384_ clknet_leaf_15_wb_clk_i net675 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_32_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08022__X _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11005_ net390 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
XANTENNA__05365__Y _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05697__B1 _01409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05290_ _00988_ _00989_ _00982_ vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09960__RESET_B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10875__551 vssd1 vssd1 vccd1 vccd1 _10875__551/HI net551 sky130_fd_sc_hd__conb_1
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06413__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08980_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__nand4_1
XFILLER_0_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07931_ _03314_ _03484_ _03485_ net256 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07862_ net277 _03414_ _03416_ net275 vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__o22a_1
X_09601_ _04677_ _04678_ vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__nor2_1
XANTENNA__06716__A3 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06813_ _02479_ _02481_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__nand2_1
X_07793_ net282 _01069_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10411__Q team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09532_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[34\]
+ net270 _04638_ _04645_ net223 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__a221o_1
X_06744_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[0\]
+ _02415_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__nand2_1
XANTENNA__06387__X _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00820_ net273 vssd1 vssd1
+ vccd1 vccd1 _04605_ sky130_fd_sc_hd__and3_4
XANTENNA__07677__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06675_ net96 _02347_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout253_A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06547__B net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08414_ net474 _03643_ _03815_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__or3b_1
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05626_ net420 _00679_ _01327_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09394_ net417 _01416_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08345_ _03631_ _03662_ _03821_ _03659_ _03629_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__o221a_1
X_05557_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\] vssd1 vssd1 vccd1
+ vccd1 _01270_ sky130_fd_sc_hd__or3_2
XFILLER_0_117_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08276_ net130 _03670_ _03754_ _03654_ vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__a31o_1
X_05488_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07227_ net257 _01655_ _02276_ _02877_ _02040_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07158_ _02060_ _02112_ _02810_ _02809_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09051__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06109_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\]
+ _01791_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__nor3_1
XFILLER_0_30_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07089_ net261 _01658_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout120 _01607_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_4
Xfanout131 net133 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_4
Xfanout142 net143 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_2
Xfanout153 net155 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout164 net165 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__buf_2
Xfanout175 net177 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
Xfanout186 _01532_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_4
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_83_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05913__Y _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07841__B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06340__A1 _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10505_ clknet_leaf_14_wb_clk_i _00373_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06192__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10859__535 vssd1 vssd1 vccd1 vccd1 _10859__535/HI net535 sky130_fd_sc_hd__conb_1
XFILLER_0_111_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10436_ clknet_leaf_44_wb_clk_i _00320_ net384 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10367_ clknet_leaf_22_wb_clk_i net677 net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10298_ clknet_leaf_39_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[11\]
+ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10231__Q team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07659__A1 _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06367__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06460_ net267 _00755_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__nor2_2
XFILLER_0_73_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05411_ net193 _01015_ _01043_ _01114_ _01123_ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__o2111a_1
X_06391_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] _00755_
+ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__nor2_2
XFILLER_0_84_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08130_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[14\]
+ _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07479__A _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05342_ net437 _00669_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08061_ net1004 net1183 net298 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05273_ _00985_ vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07012_ _02663_ _02662_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_116_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05727__A _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\] net826
+ net447 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07914_ _01689_ _03381_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__nor2_1
X_08894_ _04212_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[4\]
+ _04209_ vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__mux2_1
X_07845_ _01077_ net113 vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout370_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07776_ _00669_ _01607_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__nand2_1
X_04988_ team_07_WB.instance_to_wrap.audio vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
XANTENNA__05462__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[28\]
+ net271 net292 net222 vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__a211o_1
XFILLER_0_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06727_ _02395_ _02396_ _02399_ _01639_ _01630_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a311o_1
XANTENNA__06277__B net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_X net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07100__A_N _02726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09446_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[0\]
+ net417 _04585_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__or3b_1
X_06658_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\] net275
+ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05609_ net445 net444 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__nor2_1
X_09377_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ _04538_ _04540_ _04542_ vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__o22a_1
XFILLER_0_136_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06589_ net124 _01654_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__nor2_2
XFILLER_0_47_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08328_ _00683_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ _03804_ _03747_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06724__C _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ net488 _00727_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06580__X _02254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10221_ clknet_leaf_0_wb_clk_i _00225_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[31\]
+ sky130_fd_sc_hd__dfrtp_2
X_10971__612 vssd1 vssd1 vccd1 vccd1 _10971__612/HI net612 sky130_fd_sc_hd__conb_1
XANTENNA__06740__B _00675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07328__S _01109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ clknet_leaf_1_wb_clk_i net698 net308 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10083_ clknet_leaf_69_wb_clk_i _00141_ net349 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05924__X _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06010__B1 _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08838__B1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10985_ net626 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07813__B2 _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10457__RESET_B net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold409 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06490__X _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ clknet_leaf_53_wb_clk_i _00310_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05547__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07041__A2 _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05960_ _01574_ _01575_ net144 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__a21o_4
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_04911_ net479 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__inv_2
X_05891_ _01579_ _01581_ _01584_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__and3_2
XFILLER_0_75_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07630_ _02070_ _03120_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__or2_1
XANTENNA__06552__A1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06552__B2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07561_ net171 _02744_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__or2_2
XFILLER_0_49_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09300_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[8\]
+ _04486_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__nand2_1
X_06512_ _02120_ _02185_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07492_ net89 net119 _02191_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09231_ net231 _04438_ _04439_ net408 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06443_ _02062_ _02076_ _02092_ _02116_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06825__B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09162_ net210 _04387_ _04388_ net401 net1117 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_118_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06374_ net135 net141 net173 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_133_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08113_ net762 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[3\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__mux2_1
X_05325_ net192 _01027_ vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09093_ _04337_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout216_A _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ _03575_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[16\]
+ net456 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__mux2_1
X_05256_ _00669_ _00967_ vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__nor2_1
XANTENNA__06841__A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05187_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] _00843_ _00898_
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] vssd1 vssd1 vccd1 vccd1
+ _00900_ sky130_fd_sc_hd__a22o_1
XANTENNA__07656__B _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ clknet_leaf_41_wb_clk_i net1017 net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09871__B _01789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _00709_ _00710_ _04234_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_cleared
+ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__a31o_1
XANTENNA__06791__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06791__B2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ net439 _01389_ _02930_ _04201_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07828_ _01057_ net219 net200 _01094_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__a22o_1
X_07759_ _01078_ _01513_ _01516_ _03313_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10770_ clknet_leaf_66_wb_clk_i _00591_ net355 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09429_ _00810_ _02961_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821__497 vssd1 vssd1 vccd1 vccd1 _10821__497/HI net497 sky130_fd_sc_hd__conb_1
XFILLER_0_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07559__B1 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10204_ clknet_leaf_84_wb_clk_i _00208_ net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10135_ clknet_leaf_59_wb_clk_i team_07_WB.instance_to_wrap.team_07.defusedGen.defusedDetect
+ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.defusedGen.defusedPixel
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10066_ clknet_leaf_38_wb_clk_i _00124_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07731__B1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10968_ net609 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_39_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10899_ net565 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05110_ net1006 _00824_ _00825_ net979 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06090_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[3\] _01772_ vssd1
+ vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold206 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold217 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[46\]
+ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold228 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[6\]
+ vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05118__A_N net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05041_ _00771_ _00772_ vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold239 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[7\]
+ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11015__641 vssd1 vssd1 vccd1 vccd1 _11015__641/HI net641 sky130_fd_sc_hd__conb_1
X_08800_ net865 _04154_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06222__B1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] _04798_ _04803_
+ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__and3_1
X_06992_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[14\] _02652_
+ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07492__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[5\] team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ net236 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__mux2_1
X_05943_ net88 _01636_ _01635_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_89_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08662_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ _00707_ _04051_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__o22a_1
X_05874_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] net148
+ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__nand2_1
X_07613_ _01647_ net103 _02762_ net149 vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__a2bb2o_1
X_08593_ _03620_ _04030_ net139 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout166_A _02055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07544_ _01646_ net102 _03101_ _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07475_ net990 _00824_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout333_A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09214_ net230 net406 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06426_ _02058_ _02091_ _02099_ _01693_ _02098_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06274__C net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ net210 net400 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06357_ net274 _02030_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout121_X net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout219_X net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05308_ _00993_ _00994_ vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__nand2_4
X_06288_ _00681_ net134 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__nor2_1
X_09076_ net212 net403 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08027_ _03564_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ net393 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__mux2_1
X_05239_ _00935_ _00931_ vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_102_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09978_ clknet_leaf_0_wb_clk_i _00083_ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_18_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__05915__A _01582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ net437 net821 net244 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06449__C _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ net498 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_28_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09466__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10753_ clknet_leaf_66_wb_clk_i team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[0\]
+ net345 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10684_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[16\]
+ net354 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07577__A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07525__C_N net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10118_ clknet_leaf_27_wb_clk_i _00156_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10049_ clknet_leaf_29_wb_clk_i _00107_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05590_ net419 _00676_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__or3_2
XFILLER_0_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07104__X _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07260_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[8\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06211_ _01890_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__inv_2
X_07191_ _02834_ _02838_ _02839_ _02842_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07487__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06142_ net114 _01801_ _01803_ net91 _01822_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__a221oi_1
XANTENNA__06391__A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06073_ team_07_WB.instance_to_wrap.team_07.maze_clear_edge_detector.inter _00803_
+ _00804_ _00806_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__or4_4
XFILLER_0_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09901_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[10\] _01777_
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[11\] vssd1 vssd1 vccd1
+ vccd1 _04888_ sky130_fd_sc_hd__o21ai_1
X_05024_ net279 _00750_ vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10414__Q team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09932__A1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09832_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[8\] _04840_ vssd1
+ vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__nand2_1
X_09763_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__inv_2
X_06975_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[6\] _02641_
+ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout283_A team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__nand2_1
X_05926_ net287 net282 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__or2_2
X_09694_ _04731_ _04741_ _04743_ _04730_ net1031 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__a32o_1
X_08645_ _04060_ _04070_ _04071_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05857_ _01524_ _01533_ _01549_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__or3_2
XFILLER_0_117_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout169_X net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[15\]
+ _03617_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05788_ _00709_ net418 _01436_ _01434_ net1159 vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__a32o_1
XANTENNA__07014__X _02671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07527_ net102 _02263_ _01708_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07458_ net453 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06409_ _01687_ _01695_ _02082_ _01647_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07389_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[2\] vssd1 vssd1 vccd1
+ vccd1 _02987_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09128_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ net403 net213 _04362_ vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09059_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10782__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11021_ net391 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07336__S _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05960__A2 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05932__X _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07162__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06476__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10805_ clknet_leaf_78_wb_clk_i _00626_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05811__C net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10736_ clknet_leaf_61_wb_clk_i _00566_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05476__A1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10667_ clknet_leaf_50_wb_clk_i _00522_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_11_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07217__A2 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10598_ clknet_leaf_54_wb_clk_i _00462_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07754__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06728__B2 _02134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09390__A2 _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06003__X _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06760_ _02426_ _02431_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__nand2_1
XANTENNA__07770__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05711_ net478 _01423_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_125_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06691_ _02079_ _02362_ _02363_ _02210_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08430_ _03756_ _03898_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__xor2_1
X_05642_ _01348_ _01353_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08361_ _00730_ _03836_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05573_ _01284_ _01285_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07312_ net685 net726 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.nxt_rand_num\[2\]
+ sky130_fd_sc_hd__nor3b_1
XFILLER_0_129_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08292_ _03720_ net416 _03671_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__or3b_1
XFILLER_0_116_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07243_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ _00719_ _02892_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06833__B net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07174_ _02824_ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06125_ _01805_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__inv_2
XANTENNA__07759__A3 _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06056_ net106 net142 _01645_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout302 _00829_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_2
X_05007_ _00738_ _00739_ _00740_ _00743_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__or4_4
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout313 net316 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_4
Xfanout324 net329 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_4
Xfanout335 net338 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_2
Xfanout346 net350 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input3_A gpio_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _04827_ _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__nor2_1
Xfanout357 net389 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_2
Xfanout368 net375 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_2
Xfanout379 net380 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\] _00763_ _00780_
+ _04777_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__and4_1
X_06958_ net105 _02628_ _02626_ _02520_ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08776__A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05068__D_N team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05909_ _01583_ net122 _01602_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__a21oi_2
X_09677_ _04731_ _04730_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06889_ _02548_ _02551_ _02558_ _02559_ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__and4b_1
X_08628_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ _04047_ _04050_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[2\]
+ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__o221a_1
XFILLER_0_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07695__A2 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06296__A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08559_ _03650_ _03961_ _04009_ vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10521_ clknet_leaf_19_wb_clk_i _00389_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06655__B1 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06743__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10452_ clknet_leaf_47_wb_clk_i _00336_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10383_ clknet_leaf_15_wb_clk_i net706 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06958__A1 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_57_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ net390 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07590__A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07135__A1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05381__Y _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07686__A2 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06894__B1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05541__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[13\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10719_ clknet_leaf_62_wb_clk_i _00550_ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07749__B _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06949__A1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06413__A3 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07930_ _03446_ _03482_ _03483_ net219 _01067_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__o32a_1
XFILLER_0_48_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07861_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\] _03281_
+ _03292_ _03415_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__or4_2
XFILLER_0_138_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09600_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[7\] _04665_ _04675_
+ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__and3_1
X_06812_ _02479_ _02481_ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05385__B1 _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07792_ net299 net118 vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__xnor2_1
X_09531_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[2\] _04640_
+ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__nand2_1
X_06743_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear_detector0.pos_y\[2\]
+ net430 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__nand2_1
XANTENNA__07126__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09462_ net893 net208 _04604_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__o21a_1
XANTENNA__07677__A2 _01723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06674_ _00755_ _01582_ net117 net110 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__o31a_1
X_08413_ _03753_ _03887_ _03751_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05625_ net419 net443 _01323_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__a21o_1
X_09393_ net417 _01416_ _01477_ _04552_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__a31o_1
X_08344_ net467 _03641_ _03660_ _03761_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__o31a_1
XFILLER_0_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05556_ _01254_ _01268_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06844__A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08275_ _03750_ _03753_ _03752_ _03716_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout413_A _00706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05487_ _00688_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ _01199_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__o21ai_1
X_07226_ net171 _01744_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07157_ _02138_ net81 _02750_ _02807_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout201_X net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06108_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[2\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__or4b_1
XFILLER_0_100_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07088_ _02134_ net81 _02732_ _02741_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06039_ net172 _01715_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__nor2_2
Xfanout110 _01615_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout121 net125 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_4
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_6
XANTENNA_input6_X net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout143 _01697_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
Xfanout165 _02745_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__buf_2
XANTENNA__06168__A2 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 net177 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_8
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_4
Xfanout198 _01518_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_8
X_09729_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\] _04767_ _04766_
+ vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_2_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08937__C _01762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06738__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07668__A2 _02260_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06754__A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07569__B _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10504_ clknet_leaf_14_wb_clk_i _00372_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_59_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10435_ clknet_leaf_48_wb_clk_i _00319_ net382 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07053__B1 _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10366_ clknet_leaf_22_wb_clk_i net723 net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10297_ clknet_leaf_39_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[10\]
+ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08856__A1 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07659__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05410_ _01006_ _01012_ _01026_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__nor3_1
XFILLER_0_28_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06390_ _02053_ _02063_ _02031_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_32_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05341_ _01028_ _01034_ _01052_ _01050_ vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__o31a_1
XANTENNA__07479__B _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08060_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ _03027_ _03583_ _03584_ vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05272_ net426 net429 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__nand2_2
X_07011_ _02656_ _02669_ _02655_ vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07595__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08962_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\] net824
+ net448 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__mux2_1
X_07913_ _01691_ _03381_ _03467_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__o21a_1
X_08893_ _00708_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[3\]
+ net482 vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07347__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10422__Q team_07_WB.instance_to_wrap.team_07.DUT_maze.mazer_locator0.activate_rand_delay
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07844_ _01076_ net109 vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__nand2_1
X_07775_ net435 net116 vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout363_A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04987_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.rand_y\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
X_09514_ net918 net207 _04634_ vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__o21a_1
X_06726_ _02107_ _02154_ _02260_ _02398_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a31oi_1
XANTENNA__05462__B team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08847__A1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ net961 net208 _04592_ vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06657_ _02066_ _02329_ _02327_ _02328_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout151_X net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05608_ net443 team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\] vssd1 vssd1
+ vccd1 vccd1 _01321_ sky130_fd_sc_hd__nor2_1
X_09376_ _04541_ net226 vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__and2b_1
X_06588_ net254 _02021_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08327_ net4 _00660_ _03743_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ _00721_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__o311a_4
XFILLER_0_47_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05539_ _01243_ _01250_ _01251_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06724__D _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ net459 _03735_ _03736_ _03695_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07209_ _02858_ _02859_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08189_ net469 net471 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\] vssd1 vssd1
+ vccd1 vccd1 _03668_ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10220_ clknet_leaf_86_wb_clk_i _00224_ net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07586__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ clknet_leaf_1_wb_clk_i net720 net308 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[10\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_7_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10082_ clknet_leaf_68_wb_clk_i _00140_ net348 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_leng\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06546__C1 _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06010__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05372__B _01014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10984_ net625 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10826__502 vssd1 vssd1 vccd1 vccd1 _10826__502/HI net502 sky130_fd_sc_hd__conb_1
XFILLER_0_69_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07813__A2 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10418_ clknet_leaf_10_wb_clk_i _00309_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_74_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08204__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10349_ clknet_leaf_40_wb_clk_i _00289_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05547__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07041__A3 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10426__RESET_B net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04910_ net741 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[0\]
+ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05890_ _00716_ _01569_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__nor2_1
XANTENNA__06659__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07107__X _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06552__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07560_ _03117_ _03118_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__or2_2
XFILLER_0_49_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06511_ _01708_ _01812_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07491_ _03045_ _03047_ _03051_ _03041_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.buttonDetect
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_75_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09230_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[5\]
+ _04435_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__nand2_1
X_06442_ _02054_ _02115_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__04907__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_86 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09161_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04384_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06373_ net203 _02046_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__nand2_2
XFILLER_0_90_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08112_ net755 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[2\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05324_ net192 _01027_ vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09092_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04333_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08043_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[18\]
+ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[22\]
+ net452 vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__mux2_1
X_10994__635 vssd1 vssd1 vccd1 vccd1 _10994__635/HI net635 sky130_fd_sc_hd__conb_1
X_05255_ net437 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1
+ vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout111_A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05186_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] _00840_ _00898_
+ _00833_ vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__a22o_1
XANTENNA__07656__C _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06592__A_N _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09994_ clknet_leaf_42_wb_clk_i _00033_ net386 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10167__RESET_B net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07953__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ net973 _04237_ _04239_ vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout480_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout199_X net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ net445 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[0\] vssd1 vssd1
+ vccd1 vccd1 _04201_ sky130_fd_sc_hd__xnor2_1
X_07827_ _01095_ net189 vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__nor2_1
XANTENNA__06288__B net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ _01066_ net216 vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06709_ _02134_ _02149_ net83 _02139_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07689_ _03203_ _03221_ _03246_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.defusedGen.defusedDetect
+ sky130_fd_sc_hd__or3_1
X_09428_ _04568_ _04569_ _04578_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_137_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09359_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ _04525_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08048__A2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09548__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07559__A1 _02135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10590__RESET_B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ clknet_leaf_86_wb_clk_i _00207_ net305 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10134_ clknet_leaf_27_wb_clk_i net768 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input41_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06782__A2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ clknet_leaf_38_wb_clk_i _00123_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__07731__A1 _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10967_ net608 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_67_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10898_ net564 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_39_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10978__619 vssd1 vssd1 vccd1 vccd1 _10978__619/HI net619 sky130_fd_sc_hd__conb_1
XFILLER_0_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10678__RESET_B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08860__C _00960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07757__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold207 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold218 _00506_ vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 _00095_ vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__dlygate4sd3_1
X_05040_ _00768_ _00769_ _00770_ vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__nand3_2
XANTENNA__06470__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06470__B2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06222__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06991_ _02653_ _02654_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__nand2_1
XANTENNA__08221__X _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06773__A2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ net1096 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ net237 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__mux2_1
XANTENNA__07970__B2 _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07492__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05942_ _00755_ _01621_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__nor2_4
XANTENNA__06389__A _02060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08661_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[8\]
+ _04085_ _04087_ _04088_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__a22oi_2
X_05873_ _01562_ _01564_ _01560_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__a21o_1
XANTENNA__07183__C1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07612_ _03118_ _03153_ _03169_ _02229_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__o211a_1
X_08592_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[16\]
+ _03618_ net889 vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07543_ net128 _01701_ net165 vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06395__Y _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout159_A _01558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07474_ net484 net1169 vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ net406 _04426_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06425_ net202 _01745_ _01663_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_107_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout326_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09144_ net333 _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_20_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06356_ net280 net283 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__nand2_4
XFILLER_0_115_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05307_ _00990_ _01014_ _01019_ vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__or3_2
X_09075_ net332 _04324_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06287_ _00681_ net134 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout114_X net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08026_ _00706_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ net295 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ _03563_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05238_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ _00948_ _00949_ _00950_ vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__a311o_1
XFILLER_0_114_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05169_ _00866_ _00880_ _00881_ _00857_ vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ clknet_leaf_85_wb_clk_i _00082_ net315 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07961__A1 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07961__B2 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05915__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] net735 net244
+ vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08859_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ net297 net294 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ _04190_ vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__a221o_1
XANTENNA__07713__A1 _03256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10821_ net497 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
XANTENNA__05931__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10752_ clknet_leaf_71_wb_clk_i _00582_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10683_ clknet_leaf_64_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[15\]
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10771__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08977__A0 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10700__RESET_B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06204__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__A _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07401__B1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ clknet_leaf_28_wb_clk_i _00155_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05825__B net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10048_ clknet_leaf_28_wb_clk_i _00040_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.idle
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold90 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[7\] vssd1 vssd1
+ vccd1 vccd1 net760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06210_ net110 _01801_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__or2_1
XANTENNA__06691__A1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07768__A _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07190_ _02840_ _02841_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06141_ net114 _01801_ _01821_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07487__B _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10434__CLK clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06391__B _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06072_ net243 _01749_ _01758_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__or3_4
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09900_ net1069 net154 net151 _04887_ vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05023_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\] net284
+ vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09831_ _04840_ _04841_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\]
+ net247 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__04920__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__A1 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09762_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\]
+ _04785_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__and3_1
X_06974_ _02641_ _02642_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__nor2_1
X_08713_ _04129_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ _04128_ vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__mux2_1
X_05925_ _01616_ _01617_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__nand2_2
X_09693_ _04742_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08644_ _04070_ _04071_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__nand2_1
X_05856_ _01533_ _01549_ _01524_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08575_ _03997_ _04020_ _03996_ vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_25_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05787_ net489 _01435_ _01484_ _01433_ net490 vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_25_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07526_ _01708_ net102 vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07457_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ net396 net298 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ _03029_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[6\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06408_ net124 _01701_ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_40_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07388_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[2\] vssd1 vssd1 vccd1
+ vccd1 _02986_ sky130_fd_sc_hd__a21o_1
X_09127_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__xnor2_1
X_06339_ net188 _01741_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__nand2_2
X_09058_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[10\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[7\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__and4_1
XFILLER_0_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08009_ _03556_ _03557_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout91_A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ net391 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05926__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08302__A team_07_WB.instance_to_wrap.team_07.heartPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07147__C1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08956__B net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__B1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06757__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07162__A2 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06476__B _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10804_ clknet_leaf_78_wb_clk_i _00625_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10735_ clknet_leaf_72_wb_clk_i _00565_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07588__A _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10666_ clknet_leaf_50_wb_clk_i _00521_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09611__A1 _04666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10597_ clknet_leaf_54_wb_clk_i _00461_ net366 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06425__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10250__Q team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05710_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\] _01417_
+ _01421_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__or4_2
XFILLER_0_76_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07770__B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06690_ net88 _02148_ net253 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_125_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06667__A _02108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05571__A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05641_ _01348_ _01353_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06361__B1 _01683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08360_ _01260_ _03724_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__o21ai_1
X_05572_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\] vssd1 vssd1 vccd1
+ vccd1 _01285_ sky130_fd_sc_hd__or3b_2
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07311_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[2\]
+ _02931_ _02934_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[2\]
+ sky130_fd_sc_hd__a21o_1
X_08291_ _03759_ _03764_ _03768_ _03630_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07242_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06664__A1 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07173_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[29\] net300 _02673_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[5\]
+ _02823_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08106__B _02671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06416__A1 _02087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06124_ net117 _01797_ _01804_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06055_ net199 net205 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__nand2_4
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05006_ net32 net31 _00741_ _00742_ vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout303 net305 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_4
Xfanout314 net316 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_4
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_4
Xfanout336 net338 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_4
Xfanout347 net350 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_4
X_09814_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\]
+ _04826_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__and3_1
Xfanout358 net363 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_4
Xfanout369 net370 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_4
X_09745_ net984 _04776_ _04778_ vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout181_X net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06957_ _02497_ _02627_ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__nor2_1
XANTENNA__08776__B _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05908_ _01569_ _01578_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__xnor2_1
X_09676_ _00762_ _04710_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__nor2_2
X_06888_ net90 _02544_ _02554_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05481__A _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08627_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ _04049_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__or2_1
X_05839_ _01527_ _01530_ _00714_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08558_ _03613_ _04008_ net139 vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07509_ net169 _01739_ _02041_ _02085_ _01690_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_64_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08489_ net54 _02670_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10520_ clknet_leaf_17_wb_clk_i _00388_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10451_ clknet_leaf_47_wb_clk_i _00335_ net374 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08731__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10382_ clknet_leaf_15_wb_clk_i net671 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05359__C _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05927__Y _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout94_X net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold390 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[9\] vssd1 vssd1
+ vccd1 vccd1 net1060 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net638 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_88_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_73_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09562__S net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07590__B _02109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05697__A2 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10718_ clknet_leaf_60_wb_clk_i _00549_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08207__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10649_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[6\]
+ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10245__Q team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07860_ _03330_ _03331_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_127_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06811_ net286 _00695_ _02481_ _02480_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__a31o_1
X_07791_ _03341_ _03342_ _03343_ _03344_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__or4_2
XFILLER_0_78_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09530_ net970 net206 _04644_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__o21a_1
X_06742_ _02413_ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__inv_2
XANTENNA__06397__A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07126__A2 _00749_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09461_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[5\]
+ net272 _04603_ net290 net220 vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__a221o_1
X_06673_ _02129_ _02312_ _02329_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__or3b_1
XANTENNA__07677__A3 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05624_ net444 _01336_ _01333_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__o21ai_1
X_08412_ _00048_ _03878_ _03886_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09392_ _01415_ _01476_ net479 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08343_ net468 _03816_ _03819_ _03664_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__o22a_1
X_10843__519 vssd1 vssd1 vccd1 vccd1 _10843__519/HI net519 sky130_fd_sc_hd__conb_1
XFILLER_0_4_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10772__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05555_ _01266_ _01267_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout141_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout239_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08274_ net54 _00702_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__nor2_4
X_05486_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ _00689_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07225_ _02860_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout406_A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07156_ _02062_ _02186_ _02808_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__and3_1
X_06107_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[24\] _01787_
+ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07087_ _01618_ _02214_ _02735_ _02107_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06038_ _01668_ _01716_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_1111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout100 net101 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout111 net113 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout122 net125 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_2
XFILLER_0_100_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout133 _01577_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout144 _01649_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_4
Xfanout155 _04868_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_2
Xfanout166 _02055_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_4
XANTENNA__06168__A3 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout177 net179 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_4
Xfanout188 net189 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_4
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ _03455_ _03542_ _03543_ _03466_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_2_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09728_ _00772_ _00779_ _00783_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_83_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09511__B1 _04584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _04719_ _04718_ net1172 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08078__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ clknet_leaf_14_wb_clk_i _00371_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10898__564 vssd1 vssd1 vccd1 vccd1 _10898__564/HI net564 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_59_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09578__B1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09557__S net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10434_ clknet_3_0_0_wb_clk_i _00318_ net311 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07053__A1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10365_ clknet_leaf_22_wb_clk_i net683 net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10296_ clknet_leaf_39_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[9\]
+ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05392__Y _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07106__A _01630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08856__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10285__RESET_B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06367__D net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06945__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10946__587 vssd1 vssd1 vccd1 vccd1 _10946__587/HI net587 sky130_fd_sc_hd__conb_1
XFILLER_0_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05340_ _01052_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05271_ net426 net427 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__xor2_2
X_07010_ _02656_ _02669_ vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06680__A _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08961_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\] net812
+ net447 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07912_ net147 _03405_ _03464_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__a21oi_1
X_08892_ _04211_ net974 _04209_ vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__mux2_1
X_07843_ _03345_ _03397_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout189_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ net105 _03321_ _03326_ net106 vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__o2bb2a_1
X_04986_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09513_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[27\]
+ net271 _04584_ net224 vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a211o_1
X_06725_ _02031_ _02264_ _02397_ _02128_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_79_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08847__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06656_ _02269_ _02284_ _02286_ _02265_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__o22ai_4
X_09444_ net290 _04590_ net272 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[0\]
+ net220 vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05607_ net446 _01314_ _01315_ _01319_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__o32a_1
X_09375_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ _04538_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__and2_1
X_06587_ net254 _02021_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout144_X net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05538_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ _01108_ _00797_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__o21a_1
X_08326_ _03674_ _03802_ _03713_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08257_ _01296_ _01302_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05469_ _01042_ _01051_ _01180_ _01181_ _01032_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_132_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07208_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00829_ _00943_ _02857_
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08188_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__nor2_2
XFILLER_0_15_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06590__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07139_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] net302 net398 _02790_
+ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__a22o_1
XANTENNA__05918__B net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10241__SET_B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07586__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ clknet_leaf_3_wb_clk_i net708 net310 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[9\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05637__C team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ clknet_leaf_27_wb_clk_i _00139_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.tft_reset
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10983_ net624 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865__541 vssd1 vssd1 vccd1 vccd1 _10865__541/HI net541 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_48_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05521__B2 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10417_ clknet_leaf_12_wb_clk_i _00308_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_74_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06005__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10348_ clknet_leaf_40_wb_clk_i _00288_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06785__B1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ clknet_leaf_86_wb_clk_i _00271_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11009__639 vssd1 vssd1 vccd1 vccd1 _11009__639/HI net639 sky130_fd_sc_hd__conb_1
XFILLER_0_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06510_ _02135_ _02178_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__nor2_1
X_07490_ _02034_ _02035_ _02231_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__a31o_1
XANTENNA__06675__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06441_ _01734_ net166 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09160_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[5\]
+ _04384_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__or2_1
X_06372_ _01642_ _02045_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08111_ net771 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[1\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__mux2_1
X_05323_ _01008_ _01013_ vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09091_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[5\]
+ _04333_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08042_ _03574_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[9\]
+ net393 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05254_ net437 team_07_WB.instance_to_wrap.team_07.DUT_maze.map_select\[0\] vssd1
+ vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__nor2_2
XANTENNA__04923__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05297__Y _01010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05185_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[7\] team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout104_A _01694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ clknet_leaf_40_wb_clk_i _00032_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_122_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08944_ net973 _04237_ net491 vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06528__B1 _02060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ net439 _01389_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__nor2_1
X_07826_ net161 _03367_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__or2_1
X_04969_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\] vssd1
+ vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
X_10849__525 vssd1 vssd1 vccd1 vccd1 _10849__525/HI net525 sky130_fd_sc_hd__conb_1
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ _01077_ net183 vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__nand2_1
X_06708_ net85 _02214_ net83 net266 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07688_ _03233_ _03237_ _03240_ _03245_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__or4_1
XANTENNA__06585__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09427_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\]
+ _04577_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__and2_1
XANTENNA__10340__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06639_ _01596_ _01599_ _01603_ net115 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__or4_4
XFILLER_0_63_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09358_ net226 _04527_ _04528_ net408 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06059__A2 _01633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08309_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[2\] _03683_ vssd1
+ vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_43_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09289_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ _04475_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05929__A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10202_ clknet_leaf_84_wb_clk_i _00206_ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06767__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ clknet_leaf_27_wb_clk_i _00171_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05935__Y _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09705__B1 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ clknet_leaf_37_wb_clk_i _00122_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_input34_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05990__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07731__A2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10966_ net607 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XANTENNA__06495__A _02119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10897_ net654 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07103__B net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold208 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold219 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[17\]
+ vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06470__A2 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06006__Y _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10647__RESET_B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06222__A2 _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06990_ _01485_ _02651_ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__nand2b_1
X_05941_ net95 net93 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__nand2_4
XANTENNA__07492__C _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06389__B _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08660_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[6\]
+ _04047_ _04050_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ _04086_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__o221a_1
X_05872_ _01560_ _01565_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__nor2_2
X_07611_ _01566_ net135 _01669_ _01672_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08591_ _03607_ _04029_ net140 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07542_ net184 _02048_ _02887_ _01798_ _02743_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__o221a_1
XANTENNA__04918__A team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10961__602 vssd1 vssd1 vccd1 vccd1 _10961__602/HI net602 sky130_fd_sc_hd__conb_1
X_07473_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[0\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[2\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09212_ _04423_ _04424_ _04425_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07013__B team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.idle vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06424_ _02043_ _02096_ _02097_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__or3b_1
XFILLER_0_118_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09143_ _04372_ _04373_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06355_ _02008_ _02029_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recMOD.modHighlightDetect
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout221_A _04582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05249__B1 _00961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06446__C1 _02110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05306_ _00993_ _00994_ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__or2_2
X_09074_ _04321_ _04322_ _04323_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06286_ team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[3\] team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[4\]
+ team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[5\] vssd1 vssd1 vccd1 vccd1
+ _01962_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05237_ _00907_ _00911_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\]
+ _00686_ vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_13_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08025_ net455 net452 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout107_X net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05168_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\]
+ _00856_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\]
+ vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__a32o_1
XANTENNA__06749__B1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05099_ net482 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[9\]
+ _00821_ _00817_ net989 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__a32o_1
X_09976_ clknet_leaf_90_wb_clk_i _00081_ net307 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08927_ net1145 net263 _04233_ vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08858_ net395 net393 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__o21a_1
XANTENNA__07713__A2 _03258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07809_ net275 _03354_ _03363_ net277 vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__o22a_1
X_08789_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\] _04139_ net965
+ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10820_ net496 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
XANTENNA__09466__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07477__A1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ clknet_leaf_71_wb_clk_i _00581_ net346 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10682_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[14\]
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07577__C net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05378__B _01083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09565__S net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_wb_clk_i_X clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05394__A _01000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ clknet_leaf_27_wb_clk_i _00154_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10047_ clknet_leaf_26_wb_clk_i net754 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.cs
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold80 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[16\]
+ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[0\] vssd1
+ vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06496__Y _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07114__A _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949_ net590 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_46_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08953__A_N net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10248__Q team_07_WB.instance_to_wrap.team_07.display_num_bus\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07768__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06140_ _01806_ _01820_ _01807_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05288__B _01000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06071_ _01197_ _01240_ _01755_ _01757_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05022_ net277 _00755_ vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__nor2_1
XANTENNA__07784__A _01058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09830_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[7\] _04838_ net269
+ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10410__RESET_B net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05403__B1 _01068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09761_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] _04788_ _04789_
+ net249 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06973_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\] net266
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] vssd1 vssd1
+ vccd1 vccd1 _02642_ sky130_fd_sc_hd__a21oi_1
X_08712_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ net243 vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__nor2_1
X_05924_ _01616_ _01617_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__and2_4
X_09692_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\] _04736_ vssd1 vssd1
+ vccd1 vccd1 _04742_ sky130_fd_sc_hd__and4_1
X_08643_ _01465_ _01475_ net478 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__o21a_4
X_05855_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[9\] net186
+ net178 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] vssd1
+ vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout171_A _01681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08574_ _03617_ _04019_ net140 vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__a21oi_1
X_05786_ net486 net488 team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\] net476 vssd1
+ vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_25_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07525_ net163 _01689_ net167 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__or3b_1
XANTENNA__10937__X net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07456_ net455 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__and2b_1
XFILLER_0_92_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06407_ net126 _01702_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_40_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07387_ net951 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\] _02985_
+ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[1\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05479__A team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_cleared vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09126_ net213 _04360_ _04361_ net400 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__a32o_1
X_06338_ net184 _01742_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_92_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09057_ _04307_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07631__A1 _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06269_ _00684_ net133 _01928_ net159 _01945_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__o221a_1
XFILLER_0_124_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07694__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08008_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[6\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05926__B net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07395__B1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09959_ clknet_leaf_86_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[28\]
+ net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[28\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__07147__B1 _02761_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05942__A _00755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07698__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__B2 _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ clknet_leaf_78_wb_clk_i _00624_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10734_ clknet_leaf_72_wb_clk_i _00564_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06122__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10665_ clknet_leaf_50_wb_clk_i _00520_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_min\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_11_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ clknet_leaf_52_wb_clk_i _00460_ net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_108_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05640_ _01350_ _01351_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06361__A1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05571_ net421 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] vssd1 vssd1 vccd1
+ vccd1 _01284_ sky130_fd_sc_hd__or3b_2
XFILLER_0_59_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07310_ _02934_ _02935_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[1\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08290_ net474 net472 _03631_ _03659_ _03767_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__o32a_1
XFILLER_0_46_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08227__X _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07241_ _02871_ _02886_ _02891_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[3\]
+ sky130_fd_sc_hd__or3_1
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07172_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[37\] net302 net301 team_07_WB.instance_to_wrap.team_07.label_num_bus\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06123_ net127 _01701_ net173 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__a21o_2
XANTENNA__06416__A2 _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07613__B2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06054_ net198 net203 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__nor2_2
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05005_ net28 net29 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout304 net305 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_4
Xfanout315 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_2
Xfanout326 net328 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_4
Xfanout337 net338 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_4
X_09813_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ _04825_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[2\] vssd1 vssd1
+ vccd1 vccd1 _04829_ sky130_fd_sc_hd__a31o_1
Xfanout348 net349 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_4
Xfanout359 net363 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_2
X_09744_ _00652_ _04777_ net248 vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__o21bai_1
X_06956_ _02520_ _02619_ _02620_ _02622_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__or4b_1
XANTENNA__06858__A net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05907_ _01590_ _01598_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09675_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _01766_ _04709_
+ _04704_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__a31o_2
XANTENNA__08877__B1 _02930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06887_ _02552_ _02557_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout174_X net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ _01249_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__and2_1
XANTENNA__05481__B _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05838_ _01527_ _01530_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__nand2_2
XFILLER_0_96_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08557_ net1173 _03612_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05769_ _01467_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[7\]
+ _01462_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__or3b_1
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07508_ _02036_ _02262_ net164 vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08488_ net814 net130 _03958_ net54 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06593__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06655__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07439_ _03018_ net233 _03017_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[20\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_130_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07852__B2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10450_ clknet_leaf_47_wb_clk_i _00334_ net368 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_116_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09109_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[10\]
+ _04347_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__or2_1
X_10381_ clknet_leaf_15_wb_clk_i net710 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10900__566 vssd1 vssd1 vccd1 vccd1 _10900__566/HI net566 sky130_fd_sc_hd__conb_1
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05937__A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold380 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] vssd1 vssd1
+ vccd1 vccd1 net1050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\] vssd1 vssd1
+ vccd1 vccd1 net1061 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout87_X net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ net390 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05375__C _01014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09144__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_42_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_103_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10717_ clknet_leaf_60_wb_clk_i _00548_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10648_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[5\]
+ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06008__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10579_ clknet_leaf_60_wb_clk_i _00014_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06810_ net282 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1 vssd1
+ vccd1 vccd1 _02481_ sky130_fd_sc_hd__or2_1
X_07790_ _03341_ _03342_ _03343_ _03344_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__nor4_1
XANTENNA__06582__B2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06741_ _02411_ _02412_ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__or2_2
XANTENNA__08859__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06397__B _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07126__A3 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[3\]
+ _04585_ _04589_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__or3_1
X_06672_ _02342_ _02344_ _02327_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__a21o_1
X_08411_ net490 net464 _03715_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__o22a_1
X_05623_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[9\] _01316_
+ _01334_ _01335_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__a211o_1
X_09391_ net417 _01416_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08342_ net467 _03766_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__nand2_1
X_10882__558 vssd1 vssd1 vccd1 vccd1 _10882__558/HI net558 sky130_fd_sc_hd__conb_1
XFILLER_0_129_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05554_ _01255_ _01265_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05485_ _00688_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ _00689_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__and3_1
XANTENNA__07834__A1 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08273_ _00048_ _03751_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout134_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07224_ _02033_ _02758_ _02872_ _02874_ _02761_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__a32o_1
XFILLER_0_42_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10436__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07155_ _02134_ net81 _02741_ _02807_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07598__B1 _03144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06106_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[24\] _01787_
+ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__nor2_2
X_07086_ _01646_ net104 _02739_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06037_ net1054 _01633_ _01641_ _01727_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wireDetect\[3\]
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout101 _01600_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout112 net113 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_4
Xfanout134 net135 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_4
Xfanout145 _01566_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout156 net157 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_4
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout167 _01719_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_4
X_10817__493 vssd1 vssd1 vccd1 vccd1 _10817__493/HI net493 sky130_fd_sc_hd__conb_1
XANTENNA__10447__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 net179 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_4
X_07988_ _03376_ _03451_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__nand2_1
Xfanout189 net190 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ net248 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[0\] vssd1
+ vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__and2b_1
X_06939_ _02607_ _02609_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09658_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\] _04713_ _04714_
+ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__and3_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08609_ _01202_ _04040_ _04039_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10597__CLK clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09589_ _04669_ _04670_ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10502_ clknet_leaf_14_wb_clk_i _00370_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09027__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10433_ clknet_leaf_57_wb_clk_i _00317_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.lives\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07053__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ clknet_leaf_22_wb_clk_i net679 net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__05386__B _01000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10295_ clknet_leaf_46_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[8\]
+ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06498__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07106__B _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07513__B1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06009__Y _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05270_ net427 net429 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__nand2_2
XFILLER_0_119_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07776__B _01607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08960_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] net835
+ net448 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05864__X _01558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ _03376_ _03465_ _03464_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__a21o_1
XANTENNA__07792__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ net482 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[6\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[2\] vssd1
+ vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__and3_1
XANTENNA__07347__A3 _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ _03395_ _03396_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__nor2_1
XANTENNA__06555__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07773_ _03298_ _03302_ _03327_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__a21o_1
X_04985_ net724 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
X_09512_ net914 net209 _04633_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06724_ net258 _01714_ _01804_ _02013_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06307__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09443_ net482 _00813_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__and2_1
X_06655_ _00649_ net286 _00757_ _01625_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__o31a_1
XFILLER_0_8_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout349_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05606_ net445 net442 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__nand2_1
XANTENNA__07303__Y _02930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[13\]
+ net408 vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__and2_1
XANTENNA__10337__SET_B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06586_ net88 _02148_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__nand2_2
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08325_ _03698_ _03782_ net486 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__a21oi_1
X_05537_ _01248_ _01249_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08256_ _03677_ _03730_ _03732_ _03734_ _01382_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05468_ _01085_ _01127_ _01097_ _01055_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07207_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[22\] net301 net300 team_07_WB.instance_to_wrap.team_07.label_num_bus\[30\]
+ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__a22o_1
XANTENNA__05758__Y _01457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ _03646_ _03663_ _03665_ _03659_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__a31o_1
XANTENNA__06590__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05399_ _01055_ _01095_ vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07138_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] net301 net300 team_07_WB.instance_to_wrap.team_07.label_num_bus\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07069_ _02682_ _02707_ _02712_ _02718_ _02723_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.displayDetect
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__08798__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06794__A1 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10080_ clknet_leaf_28_wb_clk_i _00138_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_7_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_6_0_wb_clk_i_X clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06589__Y _02262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06546__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06010__A3 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06111__A _01789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08299__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ net623 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XANTENNA__05950__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09141__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10906__572 vssd1 vssd1 vccd1 vccd1 _10906__572/HI net572 sky130_fd_sc_hd__conb_1
XFILLER_0_108_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06482__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05397__A _01000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08223__A1 _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ clknet_leaf_10_wb_clk_i _00307_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_115_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10347_ clknet_leaf_45_wb_clk_i _00287_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06005__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10278_ clknet_leaf_84_wb_clk_i _00270_ net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10762__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07117__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06021__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06440_ _02087_ _02112_ _02113_ _01711_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06371_ net188 _02044_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ net786 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.data\[0\] team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spiDataSet
+ vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05322_ net431 _00991_ _01022_ _01033_ vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__a31o_1
XANTENNA__08462__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09090_ net212 _04334_ _04335_ net399 net891 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08041_ net413 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[15\]
+ net294 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__a221o_1
X_05253_ net437 net436 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__nor2_2
XFILLER_0_114_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10292__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05184_ _00894_ _00895_ _00896_ _00891_ _00887_ vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09992_ clknet_leaf_41_wb_clk_i _00031_ net381 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06776__B2 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08943_ net995 _04235_ _04238_ vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08874_ net440 _01372_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06528__A1 _01705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ _03366_ _03378_ _03376_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__or3b_2
X_07756_ _03308_ _03310_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__or2_1
X_04968_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
XANTENNA__09478__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06707_ net175 _01737_ _02013_ _02044_ net258 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__o2111a_1
X_07687_ _03242_ _03243_ _03244_ _03129_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__o31a_1
XFILLER_0_56_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06585__B _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ _04567_ _04570_ _04576_ _00705_ _04577_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__a221oi_1
X_06638_ _02303_ _02307_ _02310_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06700__A1 _01740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09357_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ _04525_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06569_ _02050_ _02090_ _02079_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08308_ net421 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\] _03785_ vssd1
+ vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_23_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09288_ net228 _04478_ _04479_ net402 net1077 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__a32o_1
XFILLER_0_117_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08239_ net476 _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__nand2_2
XFILLER_0_105_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05929__B net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10785__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ clknet_leaf_86_wb_clk_i _00205_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06767__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10132_ clknet_leaf_27_wb_clk_i _00170_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05945__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10063_ clknet_leaf_36_wb_clk_i _00121_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05990__A2 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07192__A1 _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05951__Y _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07731__A3 _01625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10965_ net606 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_35_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10896_ net653 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_39_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold209 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[40\]
+ vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08930__S net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06016__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06222__A3 _01828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05940_ net99 net89 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07707__B1 _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05293__C _01005_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05871_ _01562_ _01564_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__and2_1
XANTENNA__07183__A1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07610_ _03098_ _03144_ _03165_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__o2bb2a_1
X_08590_ net817 _03606_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07613__A1_N _01647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07541_ net184 _02048_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07472_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[35\]
+ net294 _03037_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[39\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09211_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ net3 vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__and2_1
X_06423_ net168 _02036_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__nand2_1
XANTENNA__06692__Y _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09142_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ net5 vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06354_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.mod_row _02010_ _02027_
+ _02028_ _02026_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_20_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05305_ _01007_ _01017_ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__or2_1
XANTENNA__06446__B1 _02088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09073_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ net4 vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06285_ _01611_ _01922_ _01960_ _01961_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.buttonHighlightDetect
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout214_A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08024_ net453 net451 vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__nor2_1
X_05236_ _00918_ _00923_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05167_ _00871_ _00878_ _00879_ _00864_ _00861_ vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__a32o_1
XFILLER_0_13_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05098_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[20\]
+ _00817_ _00823_ net979 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__a22o_1
X_09975_ clknet_leaf_87_wb_clk_i _00080_ net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_08926_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[2\]
+ net241 _04228_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__and3_1
X_08857_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[36\]
+ net298 net295 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[32\]
+ _04189_ vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__a221o_1
XANTENNA__10357__RESET_B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08371__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07808_ _03355_ _03356_ _03362_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__or3_2
X_08788_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\]
+ _04139_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__or3_2
X_07739_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[2\] _03292_
+ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10750_ clknet_leaf_68_wb_clk_i _00580_ net344 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07477__A2 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09409_ _04556_ _04564_ _02962_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10681_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[13\]
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06123__X _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10115_ clknet_leaf_28_wb_clk_i _00153_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10780__RESET_B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10046_ clknet_leaf_26_wb_clk_i net790 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_dc
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07165__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10098__RESET_B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold70 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[19\] vssd1 vssd1
+ vccd1 vccd1 net740 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold81 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold92 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[4\] vssd1
+ vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__dlygate4sd3_1
X_10984__625 vssd1 vssd1 vccd1 vccd1 _10984__625/HI net625 sky130_fd_sc_hd__conb_1
XANTENNA__05715__A2 _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__RESET_B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07114__B _02282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ net589 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_128_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07468__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10879_ net555 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08226__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06428__B1 _02054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06070_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[0\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.stage\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__or3b_1
XANTENNA_1 _00990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05021_ net287 net284 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__nand2_4
XFILLER_0_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07784__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07928__B1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09760_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[10\] _04785_ _00652_
+ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a21oi_1
X_06972_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[5\] team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[4\]
+ net266 vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__and3_1
X_08711_ _01759_ _04040_ _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__nand3_1
X_05923_ _01590_ _01598_ net119 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__a21oi_1
X_09691_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[4\]
+ _04736_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\] vssd1 vssd1
+ vccd1 vccd1 _04741_ sky130_fd_sc_hd__a31o_1
X_08642_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[2\]
+ _04059_ _04068_ _04069_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__a2bb2o_4
X_05854_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _01534_
+ _01546_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__and3_1
X_08573_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[13\]
+ _03615_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05785_ _01457_ _01481_ _01483_ team_07_WB.instance_to_wrap.team_07.audio_0.ss_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout164_A net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07524_ net137 _01688_ net167 vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10439__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07455_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[1\]
+ net395 net296 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[5\]
+ _03028_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[3\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout331_A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04935__Y _00675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06406_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07386_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\]
+ net479 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09125_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ _04358_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06337_ net418 net214 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout217_X net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09056_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__and3_1
XANTENNA__07092__B1 _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06268_ net150 _01929_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08007_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__xor2_1
X_05219_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[36\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00932_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06199_ _01681_ _01873_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08302__C team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ clknet_leaf_90_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[25\]
+ net306 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ sky130_fd_sc_hd__dfstp_1
X_08909_ net438 _01398_ _01403_ team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__a31o_1
X_10968__609 vssd1 vssd1 vccd1 vccd1 _10968__609/HI net609 sky130_fd_sc_hd__conb_1
XANTENNA__07147__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ _01775_ _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__nand2_1
XANTENNA__05942__B _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__A2 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10802_ clknet_leaf_78_wb_clk_i _00623_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08745__S net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07502__X _03062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10733_ clknet_leaf_78_wb_clk_i _00563_ net341 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07221__Y _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10664_ clknet_leaf_51_wb_clk_i _00519_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_125_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07607__C1 _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_88_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10595_ clknet_leaf_52_wb_clk_i _00459_ net370 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_45_wb_clk_i_X clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XANTENNA__06189__A2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10029_ _00049_ _00045_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07125__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06361__A2 _01653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05570_ _01282_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07240_ _02761_ _02878_ _02890_ _02781_ _02888_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07171_ net449 team_07_WB.instance_to_wrap.team_07.label_num_bus\[13\] net398 vssd1
+ vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06970__Y team_07_WB.instance_to_wrap.team_07.recFLAG.flagDetect vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06122_ net198 _01801_ _01802_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06053_ net218 net200 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__nand2_4
XFILLER_0_83_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05004_ net25 net24 net27 net26 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__or4_1
XFILLER_0_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 net323 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_2
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08574__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10631__RESET_B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09812_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] _04826_ _04828_
+ net247 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__o22a_1
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_2
Xfanout338 net339 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_2
Xfanout349 net350 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_4
X_09743_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[5\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\]
+ _04772_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__and3_1
X_06955_ _02614_ _02618_ _02624_ _02625_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__o211a_1
XANTENNA__07129__A1 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05906_ _01590_ _01598_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__and2_2
X_09674_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _01766_ _04709_
+ _04704_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__a31oi_1
X_06886_ net116 _02478_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08625_ _00707_ _04052_ _04048_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05837_ _01526_ _01529_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout167_X net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08556_ net146 _04007_ _03965_ vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05768_ _01466_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[22\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[23\] vssd1 vssd1 vccd1
+ vccd1 _01467_ sky130_fd_sc_hd__or3b_2
XFILLER_0_134_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07507_ net104 net167 _02036_ _02836_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__a22o_1
X_08487_ _03630_ _03957_ net130 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06593__B _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05699_ _00826_ _01411_ vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07438_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\]
+ _03014_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07369_ net477 _02963_ _02972_ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ net212 _04346_ _04348_ net399 net1014 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__a32o_1
X_10380_ clknet_leaf_11_wb_clk_i net757 net331 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09039_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[11\]
+ _04294_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05937__B net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold370 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[6\] vssd1 vssd1
+ vccd1 vccd1 net1040 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold381 team_07_WB.instance_to_wrap.team_07.label_num_bus\[6\] vssd1 vssd1 vccd1
+ vccd1 net1051 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11001_ net392 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
Xhold392 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_82_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10716_ clknet_leaf_60_wb_clk_i _00547_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_11_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ clknet_leaf_37_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[4\]
+ net362 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06008__B _01698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10578_ clknet_leaf_60_wb_clk_i _00013_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06668__A1_N net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06024__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05909__A2 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08308__B1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ _00674_ _00675_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05790__B1 _00827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06671_ _02009_ _02027_ _02170_ _02312_ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__or4_1
X_08410_ _03718_ _03884_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nor2_1
X_05622_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[12\] net446
+ net443 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__and3_1
X_09390_ _01417_ _01477_ _04550_ _02984_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08341_ _03661_ _03815_ _03817_ net468 _03667_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05553_ _01255_ _01265_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08272_ net491 team_07_WB.instance_to_wrap.team_07.lcdOutput.playButtonPixel vssd1
+ vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__nand2_2
XFILLER_0_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05484_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[3\]
+ _01196_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07223_ net160 net107 _02872_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout127_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07154_ _02793_ _02798_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07598__A1 _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06105_ _01787_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07085_ net144 _01664_ _01660_ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06270__A1 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06036_ net261 _01718_ _01721_ _01654_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__or4b_1
XANTENNA__06270__B2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08547__B1 net140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout102 net103 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10452__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[17\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout113 net114 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout124 net125 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_4
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_8
Xfanout146 _03626_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input1_A gpio_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 _01558_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_4
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_87_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07987_ _03457_ _03540_ _03541_ _01679_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__o22a_1
Xfanout179 net180 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_2
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06573__A2 _01690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06588__B _02021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09726_ _00652_ _00780_ _00766_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__o21bai_1
X_06938_ _02515_ _02519_ _02520_ net432 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09511__A2 _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ net1144 _04717_ _04718_ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__o21a_1
X_06869_ net274 _02486_ _02539_ _02537_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08608_ _01197_ _01240_ _04037_ _01755_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__or4b_2
X_09588_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\] _04667_ net1109
+ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__a21oi_1
X_08539_ net146 _03960_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__or2_2
XFILLER_0_132_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05013__A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10501_ clknet_leaf_15_wb_clk_i _00369_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05948__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ clknet_leaf_58_wb_clk_i _00316_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08235__C1 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07589__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10363_ clknet_leaf_22_wb_clk_i net704 net336 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__05667__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06261__A1 _00684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10294_ clknet_leaf_46_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[7\]
+ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06131__X _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06498__B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07513__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08710__B1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08474__C1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06680__C _02178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06788__C1 _01636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07910_ net132 net123 _03378_ _03406_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__a31o_1
XANTENNA__07792__B net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08890_ _04210_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[2\]
+ _04209_ vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__mux2_1
XANTENNA__06689__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05593__A team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ _01115_ net111 vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07347__A4 _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07772_ _01688_ _03321_ _03326_ _01679_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__o2bb2a_1
X_04984_ net710 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
XANTENNA__05880__X _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06723_ _02134_ _02380_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09511_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[26\]
+ _04591_ _04584_ net224 vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__a211o_1
XANTENNA__07016__C _02671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07504__A1 _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ net417 _01415_ _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_52_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06654_ _02272_ _02280_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__or2_2
XFILLER_0_8_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05605_ net439 _01317_ vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__xor2_1
X_09373_ net226 _04537_ _04539_ net409 net1013 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__a32o_1
X_06585_ net88 _02148_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout244_A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08324_ net769 net130 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05536_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01239_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08255_ _01293_ _03733_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__nor2_1
X_05467_ _01175_ _01177_ _01178_ _01179_ vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout411_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07206_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[6\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[14\]
+ net450 vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08186_ net471 net475 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05398_ _01000_ net191 _01004_ vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__or3_1
XANTENNA__08768__A0 team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07137_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[3\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[11\]
+ net449 vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07068_ _02710_ _02720_ _02722_ _02693_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_54_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07991__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06019_ net107 _01698_ _01708_ net204 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_7_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input4_X net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06546__A2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05008__A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ _04752_ _04753_ net1146 _04730_ vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__a2bb2o_1
X_10981_ net622 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_97_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05950__B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08319__A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07223__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06482__A1 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07703__A2_N _01737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ clknet_leaf_12_wb_clk_i _00306_ net330 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06234__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10346_ clknet_leaf_45_wb_clk_i _00286_ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[2\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__10092__Q team_07_WB.instance_to_wrap.team_07.lcdOutput.simonPixel\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10277_ clknet_leaf_73_wb_clk_i _00269_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10833__509 vssd1 vssd1 vccd1 vccd1 _10833__509/HI net509 sky130_fd_sc_hd__conb_1
XFILLER_0_104_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10952__593 vssd1 vssd1 vccd1 vccd1 _10952__593/HI net593 sky130_fd_sc_hd__conb_1
XANTENNA__08931__A0 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08928__S net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06021__B _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06370_ net175 _01698_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05321_ net193 _01010_ _01021_ vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__nor3_2
XFILLER_0_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08040_ net453 net451 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05252_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right _00963_
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down vssd1
+ vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__or4b_4
XFILLER_0_43_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05183_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[35\] _00890_ vssd1 vssd1
+ vccd1 vccd1 _00896_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09991_ clknet_leaf_42_wb_clk_i _00000_ net385 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06776__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ net491 _04237_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__nor2_1
X_10890__647 vssd1 vssd1 vccd1 vccd1 net647 _10890__647/LO sky130_fd_sc_hd__conb_1
XANTENNA__06212__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ net438 _01399_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07824_ net143 _03377_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04967_ net451 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
X_07755_ _01066_ net174 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout361_A net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06706_ _02128_ net83 _02235_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a21o_1
X_07686_ _02070_ _02278_ _02056_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09425_ _00705_ _04576_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__nor2_1
X_06637_ _01922_ _02259_ _02305_ _02309_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__o31a_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06013__A_N _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09356_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[8\]
+ _04525_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__nand2_1
X_06568_ _01647_ _01740_ _02132_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06882__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05519_ _01225_ _01227_ _01230_ _01231_ _01204_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__o32a_1
X_08307_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[1\] _01259_ vssd1
+ vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__nand2_1
X_09287_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ _04475_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_23_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06499_ _02163_ _02164_ _02169_ _02172_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08238_ team_07_WB.instance_to_wrap.team_07.lcdOutput.modHighlightPixel team_07_WB.instance_to_wrap.team_07.lcdOutput.modSquaresPixel
+ net489 vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08169_ net54 net52 _00702_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__or3_2
XFILLER_0_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10200_ clknet_leaf_84_wb_clk_i _00204_ net314 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.label_num_bus\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08602__A team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06767__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ clknet_leaf_27_wb_clk_i _00169_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05945__B net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10062_ clknet_leaf_36_wb_clk_i _00120_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10416__SET_B net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05961__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10964_ net605 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_98_887 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05025__X _00759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06152__B1 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10895_ net652 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_31_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07888__A _01078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10815__Q team_07_WB.instance_to_wrap.team_07.heartPixel vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06016__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07955__A1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ clknet_leaf_53_wb_clk_i net684 net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06032__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07707__A1 _02040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05870_ _01534_ _01563_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__xor2_1
XANTENNA__06967__A net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07183__A2 _01699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _01618_ _01623_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07471_ net413 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[33\]
+ net395 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[37\]
+ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09210_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ net3 vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__nor2_1
X_06422_ net104 net168 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06694__B2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ net5 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__or2_1
X_06353_ _00709_ net275 _02009_ _01607_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a211o_1
XFILLER_0_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05304_ _01012_ _01016_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__or2_1
XANTENNA__06446__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.debounce
+ net4 vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__or2_1
X_06284_ net86 _01634_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08023_ net492 _03561_ _00796_ vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__mux2_1
X_05235_ _00887_ _00891_ _00892_ _00893_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout207_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05166_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[18\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00879_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06749__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855__531 vssd1 vssd1 vccd1 vccd1 _10855__531/HI net531 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_90_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07946__B2 _00752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05097_ net482 _00814_ _00821_ vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__and3_2
X_09974_ clknet_leaf_86_wb_clk_i _00079_ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_08925_ net1010 net241 _04231_ _04232_ vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout197_X net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10460__Q team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_down
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ _03024_ net394 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[34\]
+ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08371__A1 _03777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07807_ _03357_ _03358_ _03360_ _03361_ _03359_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__a221o_1
X_08787_ _04145_ _04146_ net195 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05999_ net136 net129 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__nand2_4
XANTENNA__07044__Y _02699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ _03289_ _03291_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07669_ net163 _01688_ _03198_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09408_ team_07_WB.instance_to_wrap.team_07.sck_rs_enable _04563_ net414 team_07_WB.instance_to_wrap.team_07.sck_fl_enable
+ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__a211o_1
XANTENNA__06685__A1 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ clknet_leaf_63_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[12\]
+ net353 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09339_ _04514_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06117__A _01532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05021__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05956__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10114_ clknet_leaf_28_wb_clk_i _00152_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_10045_ clknet_leaf_26_wb_clk_i _00104_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.tft_sdi
+ sky130_fd_sc_hd__dfxtp_1
Xhold60 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[0\]
+ vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07165__A2 _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold71 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[0\]
+ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold82 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[14\]
+ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 _00113_ vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10947_ net588 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_27_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10878_ net554 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_39_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08226__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06428__A1 _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06027__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_2 _01689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10839__515 vssd1 vssd1 vccd1 vccd1 _10839__515/HI net515 sky130_fd_sc_hd__conb_1
X_05020_ net280 net278 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__nor2_2
XFILLER_0_10_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09393__A3 _01477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06600__A1 _01804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06971_ _00716_ net266 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__xnor2_1
X_08710_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[0\]
+ _01243_ _04035_ net243 vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a31o_1
XANTENNA__05872__Y _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05922_ _01597_ _01604_ net112 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__and3_4
X_09690_ _00699_ _04739_ _04740_ net250 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__a22oi_1
X_08641_ net457 _04067_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__nand2_1
X_05853_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[7\] _01546_
+ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08572_ _04013_ _04018_ _03996_ vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__o21a_1
X_05784_ _00792_ team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[3\] _01481_
+ _01482_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__or4_1
XFILLER_0_83_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07523_ net165 _02836_ _01678_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout157_A _01558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07454_ net453 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10926__576 vssd1 vssd1 vccd1 vccd1 _10926__576/HI net576 sky130_fd_sc_hd__conb_1
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06405_ _00635_ net284 _00749_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__and3_4
XFILLER_0_17_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07385_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[0\] net233 vssd1
+ vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[0\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout324_A net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07616__B1 _02262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06336_ net418 net176 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__xnor2_1
X_09124_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ _04358_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07092__A1 _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09055_ net877 net407 net252 _04306_ vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06267_ _01943_ _01940_ net257 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__and3b_1
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10896__653 vssd1 vssd1 vccd1 vccd1 net653 _10896__653/LO sky130_fd_sc_hd__conb_1
XFILLER_0_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08006_ _03554_ _03555_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__xnor2_1
X_05218_ _00929_ _00930_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[8\]
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[9\] vssd1 vssd1 vccd1 vccd1
+ _00931_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_102_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06224__X _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07694__C _01639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06198_ _01656_ _01829_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05149_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[4\] team_07_WB.instance_to_wrap.team_07.label_num_bus\[6\]
+ team_07_WB.instance_to_wrap.team_07.display_num_bus\[0\] vssd1 vssd1 vccd1 vccd1
+ _00862_ sky130_fd_sc_hd__mux2_1
XANTENNA__08041__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09957_ clknet_leaf_87_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[24\]
+ net304 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[24\]
+ sky130_fd_sc_hd__dfstp_1
X_08908_ net1054 _04219_ net264 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__o21a_1
X_09888_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[6\] _01774_ vssd1
+ vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nand2_1
XANTENNA__07147__A2 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ net853 _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07698__A3 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07215__B _01901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05016__A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10801_ clknet_leaf_73_wb_clk_i _00622_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10160__RESET_B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10732_ clknet_leaf_78_wb_clk_i _00562_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07231__A _02033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10663_ clknet_leaf_51_wb_clk_i _00518_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_119_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07607__B1 _02744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10594_ clknet_leaf_39_wb_clk_i _00458_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07083__A1 _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05957__Y _01651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_102_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06013__C _01696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10028_ _00048_ _00635_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_125_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07125__B _01616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10028__CLK _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08237__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07170_ _02819_ _02821_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06121_ _01800_ _01801_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06821__A1 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06052_ net216 net197 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__nor2_4
XFILLER_0_112_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05003_ net18 net17 net15 net16 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__nand4b_1
XANTENNA__08023__A0 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout306 net323 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_4
Xfanout317 net322 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_2
X_09811_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[1\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_freq\[0\]
+ _00657_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout328 net329 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_4
Xfanout339 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.nrst
+ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_4
X_09742_ net248 _04774_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__nor2_1
X_06954_ net217 _02510_ _02616_ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07129__A2 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10671__RESET_B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05905_ _01585_ _01589_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__nand2b_1
X_09673_ _04727_ _04728_ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__nor2_1
X_06885_ _02546_ _02547_ _02549_ _02555_ _02473_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout274_A _01622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08624_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[5\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[3\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[7\]
+ net457 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_85_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06888__A1 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05836_ _01521_ _01528_ _01513_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07603__X _03162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ _03612_ _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__nand2_1
X_05767_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[15\]
+ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[12\] vssd1 vssd1 vccd1
+ vccd1 _01466_ sky130_fd_sc_hd__or3b_1
XFILLER_0_77_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07506_ _01632_ _02181_ _03063_ _03064_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__o22ai_2
X_08486_ net472 _03631_ _03955_ _03956_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__o211a_1
X_05698_ _01195_ _01410_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__nand2_4
XFILLER_0_92_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07437_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[19\] team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[18\]
+ _03013_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[20\] vssd1
+ vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__a31o_1
XFILLER_0_130_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07986__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07368_ net477 _02963_ _02970_ _02973_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[1\]
+ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_131_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09107_ _04347_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__inv_2
XANTENNA__07065__A1 _01679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06319_ net198 _01977_ _01979_ _01978_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a31o_1
XANTENNA__08262__B1 _03700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07299_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[3\]
+ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[5\]
+ _01321_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__a31o_1
XANTENNA__05076__B1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09038_ net252 _04293_ _04295_ net407 net1167 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold360 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[13\] vssd1 vssd1
+ vccd1 vccd1 net1030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold382 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[12\] vssd1 vssd1
+ vccd1 vccd1 net1052 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold393 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net392 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06576__B1 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05953__B _01645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07226__A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06130__A _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07828__B1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10715_ clknet_leaf_60_wb_clk_i _00546_ net342 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10646_ clknet_leaf_41_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[3\]
+ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10577_ clknet_leaf_24_wb_clk_i _00445_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_51_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06024__B net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06567__B1 _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10429__RESET_B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08308__A1 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08859__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05790__B2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06670_ _02009_ _02313_ _02027_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__a21o_1
X_05621_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[0\] net446
+ _00679_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08340_ _03660_ _03816_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05552_ _01256_ _01264_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08271_ _03718_ _03748_ _03749_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_129_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05483_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[1\]
+ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.simon_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07222_ _01645_ _01744_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__or2_2
XFILLER_0_61_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07153_ _02802_ _02805_ _02799_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_89_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06104_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[22\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[23\]
+ _01786_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__or3_2
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ net260 net172 _02154_ _01663_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_113_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06035_ _01654_ _01719_ _01725_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout103 _01796_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout114 _01614_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_4
Xfanout125 _01595_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout136 _01576_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_8
Xfanout147 net148 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_4
XFILLER_0_129_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout158 _01558_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_87_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout169 _01707_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06221__Y _01901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07986_ net259 _03379_ _03387_ _03406_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_52_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09725_ _04733_ _04764_ vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__nor2_1
X_06937_ _02514_ _02592_ _02515_ _02513_ _02522_ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09656_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[2\] _04717_ _04716_
+ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06868_ _02536_ _02538_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__nor2_1
X_08607_ _00688_ _04037_ _04038_ _04039_ vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__o2bb2a_1
X_05819_ _00713_ _01501_ _01504_ _01512_ _01492_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__a2111o_2
X_09587_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[3\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_bm_freq\[2\]
+ _04667_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__and3_1
XANTENNA__05533__A1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06799_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] _02467_ _02469_
+ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__a21oi_2
X_08538_ net799 _03607_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08469_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[5\] _01301_ vssd1
+ vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10500_ clknet_leaf_16_wb_clk_i _00368_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10431_ clknet_leaf_58_wb_clk_i _00315_ net358 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_cleared
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05948__B net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10362_ clknet_leaf_24_wb_clk_i net717 net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06261__A2 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10293_ clknet_leaf_46_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[6\]
+ net377 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout92_X net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05964__A _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_y\[0\]
+ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05970__Y _01664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07513__A2 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05637__A_N net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05827__A2 _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10629_ clknet_leaf_49_wb_clk_i _00493_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08777__A1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06689__B net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _01050_ net118 vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__xnor2_1
XANTENNA__05593__B team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06555__A3 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ _03303_ _03324_ _03325_ _03306_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__or4b_2
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_04983_ team_07_WB.instance_to_wrap.team_07.lcdOutput.simon_light_up_state\[1\] vssd1
+ vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
X_09510_ net906 net209 _04632_ vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__o21a_1
X_06722_ _02140_ _02394_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07504__A2 _01610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_one\[2\]
+ _04549_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__and2_1
X_06653_ _02311_ _02325_ net425 net423 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a211o_1
XFILLER_0_52_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05604_ _01315_ net446 _01314_ vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__or3b_1
X_09372_ _04538_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06584_ _01618_ _02147_ _02175_ _02257_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recPLAY.playButtonDetect
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08323_ net828 _03800_ net130 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05535_ _01194_ _01247_ _01245_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout237_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08254_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wirePixel\[4\] _01304_ vssd1
+ vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__nand2_1
X_05466_ _01033_ _01052_ net436 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_31_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07205_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] net301 net300 team_07_WB.instance_to_wrap.team_07.label_num_bus\[31\]
+ _02855_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08185_ net470 net474 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__and2_1
X_05397_ _01000_ net192 _01004_ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout404_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07136_ _02730_ _02753_ _02755_ _02778_ _02789_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.memGen.labelDetect\[0\]
+ sky130_fd_sc_hd__a221o_1
XANTENNA__10463__Q team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07067_ _02689_ _02709_ _02715_ _02110_ _02721_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_54_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06018_ _01709_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06546__A3 _01665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07969_ _01113_ net186 _01681_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__o21a_1
XANTENNA__06951__B1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\] _04750_ _04731_
+ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10980_ net621 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
X_09639_ team_07_WB.instance_to_wrap.team_07.audio_0.pzl_state\[1\] _04702_ _00761_
+ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__o21a_1
XANTENNA__06703__B1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08319__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07223__B net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05024__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06482__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ clknet_leaf_12_wb_clk_i _00305_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\]
+ sky130_fd_sc_hd__dfstp_4
XTAP_TAPCELL_ROW_115_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10345_ clknet_leaf_45_wb_clk_i _00285_ net383 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.rst_cmd\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09708__B1 _04731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05442__B1 _01067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10276_ clknet_leaf_73_wb_clk_i _00268_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_10872__548 vssd1 vssd1 vccd1 vccd1 _10872__548/HI net548 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06942__B1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06021__C _01712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05320_ net193 _01025_ vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05251_ _00658_ _00794_ _00963_ vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__nor3_4
XANTENNA__07670__A1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05182_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[34\] _00886_ vssd1 vssd1
+ vccd1 vccd1 _00895_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09990_ clknet_leaf_40_wb_clk_i _00030_ net379 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08941_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[1\] team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.num_clear\[0\]
+ _04234_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ net442 net859 net246 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__mux2_1
XANTENNA__05891__X _01585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07823_ net143 _03377_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout187_A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07754_ _01066_ net178 vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__nand2_1
X_04966_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\]
+ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XANTENNA__07489__A1 _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06705_ _02013_ _02073_ _02370_ _02371_ _02377_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a41o_1
X_07685_ _01739_ _02036_ _03198_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout354_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ _04571_ _04575_ _04576_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__and3_1
X_06636_ _02108_ _02259_ _02308_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__or3b_1
XANTENNA__06161__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10458__Q team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ net1032 net412 net227 _04526_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06567_ _02051_ _02121_ _02240_ _02067_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout142_X net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08306_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_playing.playing_state\[0\] _03783_
+ _03713_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05518_ net424 _01222_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__mux2_1
X_09286_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[4\]
+ _04475_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__nand2_1
X_06498_ net204 net253 _02171_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08237_ net463 _03714_ _03715_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__or3_1
X_05449_ _01071_ _01161_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08168_ _03630_ _03648_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07119_ _02771_ _02772_ _02769_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__a21oi_4
X_08099_ net1008 net232 _03595_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[14\]
+ vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10130_ clknet_leaf_29_wb_clk_i _00168_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10061_ clknet_leaf_37_wb_clk_i _00119_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05019__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09954__SET_B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05961__B _01654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10963_ net604 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XFILLER_0_35_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08209__A_N net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10894_ net651 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07888__B net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07652__A1 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ clknet_leaf_53_wb_clk_i net725 net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[2\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__06313__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10259_ clknet_leaf_74_wb_clk_i _00251_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06032__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07470_ net1085 net295 _03036_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[38\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06421_ _02063_ _02094_ _02080_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06694__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[13\]
+ _04371_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[16\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06352_ net98 _01616_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__and2_2
Xclkbuf_leaf_6_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05303_ _01013_ _01015_ net193 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06446__A2 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07643__A1 _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06283_ net87 net276 _01957_ _01959_ net98 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a2111oi_2
X_09071_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[13\]
+ _04320_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[16\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_112_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[3\]
+ team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[1\] vssd1 vssd1
+ vccd1 vccd1 _03561_ sky130_fd_sc_hd__or2_2
X_05234_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\] net302 _00830_ vssd1
+ vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09396__A1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05165_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[19\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout102_A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05096_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00819_ vssd1 vssd1 vccd1
+ vccd1 _00822_ sky130_fd_sc_hd__nand2_1
X_09973_ clknet_leaf_84_wb_clk_i _00078_ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[12\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_90_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06223__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08924_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.rand_start_pos_x\[1\]
+ _04228_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08855_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[25\]
+ net395 net294 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[31\]
+ _04188_ vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07806_ _01048_ net116 vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08786_ net1057 _04139_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__nand2_1
X_05998_ net131 net123 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_49_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _03289_ _03291_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__nor2_1
X_04949_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ _02081_ _02260_ _02277_ _01729_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__a22o_1
XANTENNA__06134__A1 _01812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06893__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09407_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\]
+ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[5\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\]
+ _00818_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_45_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06619_ _01812_ _02283_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06685__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07599_ _03139_ _03141_ _03157_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09338_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[0\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[2\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[1\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07634__A1 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09269_ _04419_ _04429_ _04465_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__or3b_1
XFILLER_0_8_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05021__B net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08613__A _00964_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05956__B net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07398__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10113_ clknet_leaf_28_wb_clk_i _00151_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input32_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05972__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07516__X _03075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _00064_ _00642_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[16\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_76_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold50 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.r_LFSR\[9\]
+ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.debounce
+ vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07165__A3 _02758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05691__B _00796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold72 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.debounce
+ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.internalSck vssd1 vssd1
+ vccd1 vccd1 net753 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_69_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold94 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[9\]
+ vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10946_ net587 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_27_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10877_ net553 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05716__B_N _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07625__A1 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06428__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08822__B1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921__666 vssd1 vssd1 vccd1 vccd1 net666 _10921__666/LO sky130_fd_sc_hd__conb_1
XFILLER_0_26_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_3 _03069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10878__554 vssd1 vssd1 vccd1 vccd1 _10878__554/HI net554 sky130_fd_sc_hd__conb_1
XFILLER_0_22_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06600__A2 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06970_ _02570_ _02583_ _02601_ _02640_ _02572_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.recFLAG.flagDetect
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__05882__A _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05921_ _01583_ net123 _01613_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__a21o_1
X_08640_ net457 _04067_ _04066_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__o21ai_1
X_05852_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] net179
+ _01545_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09073__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08571_ _03616_ _04017_ net139 vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__a21oi_1
X_05783_ _00777_ team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[0\] team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[1\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.nxt_cnt_s_leng\[8\] vssd1 vssd1 vccd1
+ vccd1 _01482_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07522_ _02785_ _03080_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07453_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[0\]
+ net396 net297 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[4\]
+ _03025_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[2\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06404_ _02068_ _02077_ _02066_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__o21a_1
X_07384_ net414 _01475_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05122__A team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09123_ net213 _04357_ _04359_ net400 net1124 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07616__A1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06335_ net87 _02009_ net101 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07616__B2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout317_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09054_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[15\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[14\]
+ _04301_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonUp.r_counter\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__a31o_1
X_06266_ _01924_ _01925_ _01932_ _01942_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_92_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08433__A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08005_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[11\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05217_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[38\] _00863_ vssd1 vssd1
+ vccd1 vccd1 _00930_ sky130_fd_sc_hd__xnor2_1
X_06197_ _01659_ _01877_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout105_X net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08041__A1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05148_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[23\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00861_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09956_ clknet_leaf_87_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[7\]
+ net303 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_05079_ _00803_ _00804_ _00806_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_clear
+ sky130_fd_sc_hd__nor3_1
X_08907_ _01397_ _01405_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__nor2_1
X_09887_ net849 net153 net151 _04879_ vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08838_ _04178_ _04179_ net196 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08769_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[3\] net856 net245 vssd1
+ vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__mux2_1
X_10800_ clknet_leaf_73_wb_clk_i _00621_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05016__B net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10731_ clknet_leaf_79_wb_clk_i _00561_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07855__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07231__B _02775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10662_ clknet_leaf_52_wb_clk_i _00517_ net369 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.cnt_sec_ten\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_81_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07607__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10593_ clknet_leaf_39_wb_clk_i _00457_ net376 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05967__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08032__A1 _00706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990__631 vssd1 vssd1 vccd1 vccd1 _10990__631/HI net631 sky130_fd_sc_hd__conb_1
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
XANTENNA__06043__B1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XANTENNA__07240__C1 _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06013__D _01705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10027_ clknet_leaf_59_wb_clk_i _00004_ net343 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06310__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10929_ net579 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06120_ net172 net102 _01798_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_83_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06051_ _01678_ net143 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__nand2_2
XFILLER_0_112_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06044__Y _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05002_ net21 net20 net23 net22 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08023__A1 _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout307 net323 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_4
X_09810_ team_07_WB.instance_to_wrap.team_07.audio_0.error_state\[1\] net247 vssd1
+ vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__nor2_1
Xfanout318 net322 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_4
Xfanout329 net330 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07782__B1 _02191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ _04767_ _04774_ _04775_ net248 net1098 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__a32o_1
X_06953_ _02621_ _02622_ _02623_ _02619_ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a31o_1
X_05904_ _01585_ net122 _01589_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__a21o_2
XFILLER_0_119_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09672_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[8\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[7\]
+ _04725_ _04716_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a31o_1
X_06884_ _02551_ _02552_ _02554_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07534__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08623_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.light_cnt\[0\]
+ net457 vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_90_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05835_ _01521_ _01528_ _01513_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_85_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08554_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[7\]
+ _03611_ net1149 vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__o21ai_1
X_05766_ _01461_ _01462_ _01463_ _01464_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__and4b_1
XANTENNA__04956__A team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07505_ _01619_ _01922_ _02217_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_18_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08485_ _03667_ _03953_ _03925_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05697_ _00687_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_cleared _01252_
+ _01409_ _00962_ vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__o311a_1
XFILLER_0_64_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07436_ net972 _03014_ _03016_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.nxt_cnt\[19\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07367_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[1\] team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09106_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[8\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[9\]
+ _04342_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__and3_1
X_06318_ _01964_ _01971_ _01970_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07065__A2 _01904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07298_ _02926_ _02927_ _01321_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[3\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05076__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09037_ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__inv_2
X_10974__615 vssd1 vssd1 vccd1 vccd1 _10974__615/HI net615 sky130_fd_sc_hd__conb_1
XFILLER_0_14_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06249_ team_07_WB.instance_to_wrap.team_07.memGen.mem_pos\[0\] net458 vssd1 vssd1
+ vccd1 vccd1 _01926_ sky130_fd_sc_hd__or2_2
XFILLER_0_102_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold350 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_leng\[5\] vssd1 vssd1 vccd1
+ vccd1 net1020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[5\] vssd1 vssd1
+ vccd1 vccd1 net1031 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold372 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_e_leng\[6\] vssd1 vssd1 vccd1
+ vccd1 net1042 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold383 team_07_WB.instance_to_wrap.team_07.wireGen.wire_status\[1\] vssd1 vssd1
+ vccd1 vccd1 net1053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06576__A1 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06411__A net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ net465 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
XANTENNA__07226__B _01744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05027__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07828__A1 _01057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07828__B2 _01094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10714_ clknet_leaf_62_wb_clk_i _00545_ net351 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_leng\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08772__S net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10645_ clknet_leaf_41_wb_clk_i team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[2\]
+ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10576_ clknet_leaf_24_wb_clk_i _00444_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05984__X _01677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10765__CLK clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_20_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06319__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05790__A2 _00797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10469__RESET_B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05620_ team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[15\] _01316_
+ _01332_ _00679_ _00680_ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05551_ _01262_ _01263_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08270_ _00048_ _03715_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__or2_1
X_05482_ _01194_ _01192_ _01190_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__or3b_2
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07221_ _01645_ _01744_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07152_ net107 _01710_ _02767_ _02804_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a31o_1
XFILLER_0_82_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06103_ team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[20\] team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[21\]
+ _01784_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__or3_1
XFILLER_0_112_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07083_ _02065_ net81 _02732_ _02736_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06034_ net202 _01723_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08711__A _01759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout104 _01694_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06558__A1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout115 net117 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout126 net128 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06502__Y _02176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 net138 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_4
Xfanout148 net149 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_4
X_07985_ _03374_ _03539_ _03460_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__o21a_1
Xfanout159 _01558_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout384_A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[15\] net250 _04761_
+ _04763_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_52_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06936_ _02521_ _02592_ _02595_ _02606_ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__or4_1
XANTENNA__07507__B1 _02036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09655_ _04703_ _04710_ _04714_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06867_ net282 _02474_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout172_X net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _00688_ _01242_ _01755_ _04037_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__a31o_1
X_05818_ _00712_ _01496_ _01510_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__or3_1
X_09586_ net1090 _04667_ vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__xor2_1
XANTENNA__05533__A2 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_right
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06798_ _00696_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[2\] vssd1 vssd1
+ vccd1 vccd1 _02469_ sky130_fd_sc_hd__and2_1
XANTENNA__07062__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08537_ _03994_ _03993_ net985 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05749_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[12\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[11\]
+ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[10\] vssd1 vssd1 vccd1
+ vccd1 _01448_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08468_ net459 _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__or2_1
XANTENNA__06494__B1 _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07419_ team_07_WB.instance_to_wrap.team_07.timer_sec_divider_0.cnt\[13\] _03004_
+ net478 vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08399_ net487 _03873_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10430_ clknet_leaf_55_wb_clk_i _00314_ net361 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_cleared
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06406__A _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10361_ clknet_leaf_22_wb_clk_i _00038_ net339 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06261__A3 _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10292_ clknet_leaf_45_wb_clk_i team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.nxt_wire_color_bus\[5\]
+ net378 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.rand_wire_color_bus\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold180 team_07_WB.instance_to_wrap.team_07.audio_0.count_bm_delay\[11\] vssd1 vssd1
+ vccd1 vccd1 net850 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05964__B net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[5\]
+ vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06412__Y _02086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07513__A3 _02332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06721__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05698__Y _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10628_ clknet_leaf_49_wb_clk_i _00492_ net372 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.reg_data\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10559_ clknet_leaf_19_wb_clk_i _00427_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonSelect.r_counter\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06788__A1 _01626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05874__B net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06689__C net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06051__A _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ net299 net180 vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__xnor2_1
X_04982_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.random_gen_simon_0.nxt_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
X_06721_ net177 _01702_ _02014_ _02393_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09440_ net917 net220 net290 _04588_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__a22o_1
X_06652_ _02129_ _02287_ _02312_ _02319_ _02324_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__o311a_1
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05603_ net445 _00679_ vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__nor2_1
X_09371_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[12\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonBack.r_counter\[11\]
+ _04533_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__and3_1
X_06583_ net85 _02179_ _02206_ _02239_ _02256_ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_59_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08322_ _03753_ _03799_ _03769_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05534_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_up
+ _00793_ _00794_ _01231_ _01246_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08265__X _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08253_ net461 _03731_ net460 vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_31_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05465_ _00982_ _01074_ _01091_ _01073_ vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_31_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout132_A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07204_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] net302 net398 _02854_
+ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a22o_1
X_08184_ net469 net470 _03662_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06226__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05396_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ _01108_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__nor3b_4
X_07135_ _01646_ _02783_ _02784_ _02754_ _02788_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06779__A1 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07066_ net121 _01676_ net168 _02716_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__and4_1
XFILLER_0_112_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06017_ net160 net168 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_54_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10310__CLK clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06400__B1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08940__A2 _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07968_ _01113_ net178 _03371_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__a21o_1
X_09707_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[9\] team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[10\]
+ _04749_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__and3_1
X_06919_ _02576_ _02577_ _02589_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__o21ba_1
X_07899_ _03383_ _03386_ _03453_ _03452_ _03387_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__o32a_1
XFILLER_0_69_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09638_ _00654_ _00764_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__and2_1
XANTENNA__06703__B2 _02079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09569_ _04612_ _04626_ _04657_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07223__C _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_wb_clk_i_X clknet_leaf_54_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10413_ clknet_leaf_12_wb_clk_i _00304_ net328 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_y\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05975__A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ clknet_leaf_54_wb_clk_i _00284_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wireGen.wire_pos\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10275_ clknet_leaf_73_wb_clk_i _00267_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout490 net491 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_2
XFILLER_0_75_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08695__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08447__A1 _03630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06972__C net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05250_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_left
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_select team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.reg_edge_back
+ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__or3_2
XFILLER_0_43_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08960__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07670__A2 _02277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06046__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05181_ _00892_ _00893_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08940_ net1097 _04234_ _04236_ vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__o21a_1
XANTENNA__06052__Y _01741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08871_ net444 net818 net245 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__mux2_1
X_07822_ _01095_ net158 vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07753_ _01067_ _01543_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__nor2_1
X_04965_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.initSeqCounter\[4\] vssd1
+ vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
X_06704_ _02271_ _02373_ _02374_ _02376_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__and4_1
X_07684_ _03131_ _03172_ _03241_ _03126_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__o31a_1
XANTENNA__07489__A2 _02082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09423_ _00808_ _04567_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06635_ _02266_ _02293_ _02300_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_17_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout347_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09354_ _04524_ _04525_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__nor2_1
X_06566_ net204 _02124_ _02194_ _02097_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08305_ net486 _03776_ _03781_ _03770_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__o31a_1
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05517_ _01204_ _01229_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09285_ net228 _04476_ _04477_ net401 net949 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__a32o_1
XANTENNA__07646__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06497_ _01646_ _01734_ _01660_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout135_X net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08236_ net415 _03561_ net490 vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__a21o_1
X_05448_ _01104_ _01107_ _01100_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08870__S net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05672__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08167_ net54 net52 net53 _03627_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__o31a_1
XANTENNA__04970__Y _00709_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05379_ _00970_ _01058_ vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07118_ net278 _02106_ net82 vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__or3b_1
X_08098_ _03601_ team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.cln_cmd\[14\]
+ net232 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06621__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07049_ _01921_ _02258_ net83 net265 vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10060_ clknet_leaf_28_wb_clk_i _00118_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataDc
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__05019__B _00752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06924__A1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10962_ net603 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XANTENNA__06137__C1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[0\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10893_ net650 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_67_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06152__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07521__Y _03080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07652__A2 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ clknet_leaf_51_wb_clk_i net741 net365 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.r_LFSR\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_130_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ clknet_leaf_75_wb_clk_i _00250_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_10189_ clknet_leaf_82_wb_clk_i net713 net320 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.display_num_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07340__A1 _01175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07340__B2 _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06420_ _02084_ _02093_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06351_ net261 _02017_ _02024_ _02025_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06047__Y _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05302_ _00996_ _01014_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_20_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[11\]
+ _04319_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonDown.r_counter\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06282_ net121 _01958_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08021_ team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[2\]
+ _03560_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_num_gen.nxt_wire_num\[1\]
+ sky130_fd_sc_hd__nand2_1
XANTENNA__05654__A1 team_07_WB.instance_to_wrap.team_07.lcdOutput.wire_color_bus\[16\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05233_ _00939_ _00940_ _00945_ _00834_ _00832_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__a32o_1
X_05164_ _00854_ _00875_ _00876_ _00847_ _00845_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__a32o_1
XANTENNA__10665__RESET_B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06504__A _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05095_ team_07_WB.instance_to_wrap.team_07.sck_fl_enable _00819_ vssd1 vssd1 vccd1
+ vccd1 _00821_ sky130_fd_sc_hd__and2_1
X_09972_ clknet_leaf_83_wb_clk_i _00077_ net318 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06666__A1_N net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.start_pos_x\[0\]
+ net241 _04229_ _04231_ vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__o22a_1
XANTENNA__07159__A1 _02065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout297_A _03026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[29\]
+ net296 net393 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[27\]
+ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07564__D1 _01646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07805_ _01049_ net118 vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__nand2_1
X_08785_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[2\] _04139_ vssd1
+ vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05997_ net138 net170 _01688_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout464_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ net285 _01105_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_04948_ team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_press_detector.num_pressed\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07667_ _03065_ _03223_ _03224_ _03095_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__a22o_1
XANTENNA__07331__A1 _00965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09406_ net858 _04562_ _04558_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06618_ _02129_ _02281_ _02287_ _02067_ _02290_ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__o221a_1
XFILLER_0_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07598_ _03098_ _03143_ _03144_ _03148_ _03156_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__o221a_1
XFILLER_0_137_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09337_ net227 _04512_ _04513_ net411 net1175 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__a32o_1
XFILLER_0_30_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06549_ _00758_ _01610_ net100 vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07501__C _02009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09268_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[14\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonRight.r_counter\[12\]
+ _04418_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05302__B _01014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07634__A2 _02056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08219_ net416 _03697_ net488 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09199_ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[9\]
+ team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.r_counter\[8\]
+ _04378_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__or3_1
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10112_ clknet_leaf_28_wb_clk_i _00150_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10043_ _00063_ _00641_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__05972__B net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.dest_pos_gen.r_LFSR\[2\]
+ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_sequence_gen_0.rand_simon_sequence_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_07_WB.instance_to_wrap.team_07.DUT_button_edge_detector.buttonLeft.debounce
+ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold73 team_07_WB.instance_to_wrap.team_07.wire_game_0.wire_wire_gen_0.wire_color_gen.r_LFSR\[11\]
+ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 _00106_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.spi.dataShift\[2\] vssd1
+ vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08775__S net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10945_ net586 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_27_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_45_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06530__C1 _02164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ net552 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__07873__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05884__A1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06308__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05987__X _01680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_4 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08050__A2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05920_ _01583_ net123 _01613_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__a21oi_2
XANTENNA__05882__B _01575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__A2 net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05851_ team_07_WB.instance_to_wrap.team_07.lcdOutput.framebufferIndex\[8\] _01536_
+ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__nor2_1
X_08570_ team_07_WB.instance_to_wrap.team_07.lcdOutput.tft.remainingDelayTicks\[13\]
+ _03615_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__nand2_1
X_05782_ _01477_ _01479_ _01457_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__or3b_1
X_07521_ _01655_ net170 vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__nand2_2
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07452_ net296 vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06403_ _02074_ _02076_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07383_ _02965_ _02983_ vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.nxt_cnt\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ _04358_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__inv_2
XANTENNA__05122__B team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06334_ _00751_ net276 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__or2_4
XANTENNA__07616__A2 _01676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05627__B2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09053_ net1129 net407 net251 _04305_ vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06265_ net217 _01926_ _01930_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08004_ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[4\]
+ team_07_WB.instance_to_wrap.team_07.DUT_maze.maze_pos_gen_0.map_select_gen.r_LFSR\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__xor2_1
XANTENNA__08433__B _03857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05216_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[39\] _00860_ vssd1 vssd1
+ vccd1 vccd1 _00929_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold510 team_07_WB.instance_to_wrap.team_07.timer_ssdec_sck_divider_0.cnt\[6\] vssd1
+ vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06196_ net214 _01656_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05147_ team_07_WB.instance_to_wrap.team_07.label_num_bus\[3\] _00859_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__mux2_4
XFILLER_0_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09955_ clknet_leaf_84_wb_clk_i team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.nxt_label_num_bus\[6\]
+ net313 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.mem_game_0.mem_num_gen_0.mem_num_gen.label_num_bus\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05078_ _00672_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[0\] _00696_
+ net430 _00805_ vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__a221o_1
X_08906_ _00682_ _04218_ net245 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__a21oi_1
X_09886_ _01774_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08837_ team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[20\] team_07_WB.instance_to_wrap.team_07.audio_0.count_ss_delay\[19\]
+ _04142_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__or3_1
XANTENNA__07552__A1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08768_ team_07_WB.instance_to_wrap.team_07.display_num_bus\[2\] net798 net245 vssd1
+ vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07719_ _01065_ _01590_ _01598_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _01240_ _04064_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ clknet_leaf_79_wb_clk_i _00560_ net340 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.audio_0.cnt_pzl_freq\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10661_ clknet_leaf_2_wb_clk_i _00516_ net312 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.simon_game_0.simon_light_control_0.simon_sequence_bus\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07231__C _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06128__B net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10587__RESET_B net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10592_ clknet_leaf_40_wb_clk_i _00456_ net380 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.timer_ssdec_spi_master_0.sck_sent\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07607__A2 _02073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05967__B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XANTENNA__05983__A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06043__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XANTENNA__09517__C1 _04582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10026_ clknet_leaf_53_wb_clk_i _00003_ net364 vssd1 vssd1 vccd1 vccd1 team_07_WB.instance_to_wrap.team_07.DUT_fsm_game_control.game_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10928_ net578 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
X_10845__521 vssd1 vssd1 vccd1 vccd1 _10845__521/HI net521 sky130_fd_sc_hd__conb_1
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10859_ net535 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XANTENNA__09048__B2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06050_ _01679_ _01698_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__nor2_4
XANTENNA__06054__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_05001_ _00734_ _00735_ _00736_ _00737_ vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout308 net310 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_4
Xfanout319 net322 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_2
XFILLER_0_10_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07782__A1 _01105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ team_07_WB.instance_to_wrap.team_07.audio_0.cnt_s_freq\[4\] _04772_ vssd1
+ vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__or2_1
X_06952_ net160 _02504_ team_07_WB.instance_to_wrap.team_07.DUT_maze.dest_x\[1\] vssd1
+ vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__or3b_1
.ends

