* NGSPICE file created from team_04.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

.subckt team_04 ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14] ADR_O[15]
+ ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22] ADR_O[23]
+ ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30] ADR_O[31]
+ ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0] DAT_I[10]
+ DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17] DAT_I[18]
+ DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25] DAT_I[26]
+ DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4] DAT_I[5]
+ DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12] DAT_O[13]
+ DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20] DAT_O[21]
+ DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28] DAT_O[29]
+ DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7] DAT_O[8]
+ DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O clk en gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5]
+ gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9] gpio_oeb[0] gpio_oeb[10] gpio_oeb[11]
+ gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15] gpio_oeb[16] gpio_oeb[17] gpio_oeb[18]
+ gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21] gpio_oeb[22] gpio_oeb[23] gpio_oeb[24]
+ gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28] gpio_oeb[29] gpio_oeb[2] gpio_oeb[30]
+ gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7]
+ gpio_out[8] gpio_out[9] mem_adr_start[0] mem_adr_start[10] mem_adr_start[11] mem_adr_start[12]
+ mem_adr_start[13] mem_adr_start[14] mem_adr_start[15] mem_adr_start[16] mem_adr_start[17]
+ mem_adr_start[18] mem_adr_start[19] mem_adr_start[1] mem_adr_start[20] mem_adr_start[21]
+ mem_adr_start[22] mem_adr_start[23] mem_adr_start[24] mem_adr_start[25] mem_adr_start[26]
+ mem_adr_start[27] mem_adr_start[28] mem_adr_start[29] mem_adr_start[2] mem_adr_start[30]
+ mem_adr_start[31] mem_adr_start[3] mem_adr_start[4] mem_adr_start[5] mem_adr_start[6]
+ mem_adr_start[7] mem_adr_start[8] mem_adr_start[9] memory_size[0] memory_size[10]
+ memory_size[11] memory_size[12] memory_size[13] memory_size[14] memory_size[15]
+ memory_size[16] memory_size[17] memory_size[18] memory_size[19] memory_size[1] memory_size[20]
+ memory_size[21] memory_size[22] memory_size[23] memory_size[24] memory_size[25]
+ memory_size[26] memory_size[27] memory_size[28] memory_size[29] memory_size[2] memory_size[30]
+ memory_size[31] memory_size[3] memory_size[4] memory_size[5] memory_size[6] memory_size[7]
+ memory_size[8] memory_size[9] nrst vccd1 vssd1
XFILLER_0_118_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06883_ final_design.cpu.reg_window\[211\] final_design.cpu.reg_window\[243\] net908
+ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__mux2_1
X_09671_ net263 _04582_ _04587_ _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__and4_1
XFILLER_0_158_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10023__B _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11834__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ net605 _03257_ _03232_ _02156_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__o211a_1
XANTENNA__06928__S net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ final_design.cpu.reg_window\[897\] final_design.cpu.reg_window\[929\] net854
+ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07504_ _02002_ _02032_ _02449_ _02454_ _02453_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__o41ai_2
XTAP_TAPCELL_ROW_46_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08484_ final_design.cpu.reg_window\[131\] final_design.cpu.reg_window\[163\] net864
+ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__mux2_1
XANTENNA__12291__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07435_ final_design.cpu.reg_window\[513\] final_design.cpu.reg_window\[545\] net932
+ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10841__B2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1071_A final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout427_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1169_A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07366_ _02313_ _02314_ _02315_ _02316_ net784 net805 vssd1 vssd1 vccd1 vccd1 _02317_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_135_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06663__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07288__A1_N net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09105_ _04026_ _01367_ net260 vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__mux2_1
XANTENNA__12594__B2 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09259__B net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07297_ net767 _02247_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09036_ final_design.CPU_instr_adr\[11\] _03966_ net1049 vssd1 vssd1 vccd1 vccd1
+ _00222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout796_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold340 final_design.cpu.reg_window\[570\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10357__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 final_design.cpu.reg_window\[984\] vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_X net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold362 final_design.cpu.reg_window\[170\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 final_design.cpu.reg_window\[968\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09275__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold384 final_design.cpu.reg_window\[463\] vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 final_design.cpu.reg_window\[71\] vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 net829 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_2
Xfanout831 net835 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_4
X_09938_ _04222_ _04581_ _04586_ _04727_ _04856_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__o221a_1
Xfanout842 net845 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_4
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_2
Xfanout864 net877 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__buf_2
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_2
XFILLER_0_99_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09514__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout886 net887 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__buf_2
X_09869_ _04770_ _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__xor2_1
Xfanout897 _01437_ vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_2
Xhold1040 final_design.cpu.reg_window\[615\] vssd1 vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11321__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11744__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 final_design.cpu.reg_window\[439\] vssd1 vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 final_design.cpu.reg_window\[813\] vssd1 vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ net206 net2134 net274 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12880_ clknet_leaf_79_clk _00118_ net1249 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[14\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold1073 final_design.cpu.reg_window\[830\] vssd1 vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08619__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1084 final_design.cpu.reg_window\[112\] vssd1 vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 final_design.cpu.reg_window\[546\] vssd1 vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ net198 net2217 net268 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07289__A0 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12282__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ net187 net2045 net418 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ clknet_leaf_12_clk _00732_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[489\]
+ sky130_fd_sc_hd__dfrtp_1
X_10713_ final_design.CPU_instr_adr\[13\] _05451_ net1066 vssd1 vssd1 vccd1 vccd1
+ _05452_ sky130_fd_sc_hd__mux2_1
XANTENNA__10832__B2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11693_ net214 net636 vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input92_A memory_size[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13432_ clknet_leaf_138_clk _00663_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[420\]
+ sky130_fd_sc_hd__dfrtp_1
X_10644_ _05347_ _05385_ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11699__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12872__Q final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11388__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12585__B2 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10575_ final_design.CPU_instr_adr\[6\] _04002_ net1072 vssd1 vssd1 vccd1 vccd1 _05321_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13363_ clknet_leaf_30_clk _00594_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[351\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09169__B _03649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12314_ net1987 net204 net364 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13294_ clknet_leaf_113_clk _00525_ net1212 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[282\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12245_ net569 _06175_ net506 net372 net1472 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__a32o_1
XFILLER_0_107_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12176_ net1623 net211 net381 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__mux2_1
XANTENNA__08961__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _01487_ net665 net1030 vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__a21o_1
X_11058_ net89 net1058 vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__and2_1
XANTENNA__11848__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10009_ _04085_ _04685_ _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_153_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12273__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07220_ net759 _02164_ net754 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__o21a_1
XANTENNA__07579__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07151_ final_design.cpu.reg_window\[458\] final_design.cpu.reg_window\[490\] net936
+ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08244__A2 _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07082_ _02026_ _02031_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12328__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11829__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09744__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08203__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11551__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07984_ _02932_ _02933_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__nor2_2
XFILLER_0_38_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09382__X _04301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09723_ net551 net549 net548 net547 net453 net462 vssd1 vssd1 vccd1 vccd1 _04642_
+ sky130_fd_sc_hd__mux4_1
X_06935_ final_design.cpu.reg_window\[401\] final_design.cpu.reg_window\[433\] net919
+ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout377_A _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09654_ _04189_ _04572_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_87_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06866_ net1053 net1006 net1003 _01380_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__a31o_1
XANTENNA__06658__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08605_ _02390_ _03519_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_26_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06797_ _01744_ _01745_ _01746_ _01747_ net774 net795 vssd1 vssd1 vccd1 vccd1 _01748_
+ sky130_fd_sc_hd__mux4_1
X_09585_ _03199_ _03229_ _04503_ _04140_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__a31o_1
XFILLER_0_167_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout544_A _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11067__A1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08536_ net612 _03481_ _03483_ net532 vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__o211a_1
XANTENNA__07366__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ net625 _03415_ _03416_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12395__S net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12016__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07418_ _02365_ _02366_ _02367_ _02368_ net779 net799 vssd1 vssd1 vccd1 vccd1 _02369_
+ sky130_fd_sc_hd__mux4_1
X_08398_ final_design.cpu.reg_window\[518\] final_design.cpu.reg_window\[550\] net830
+ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire528 _03513_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07349_ _02298_ _02299_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14200__1269 vssd1 vssd1 vccd1 vccd1 _14200__1269/HI net1269 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_150_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10360_ net33 net1036 net1019 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1
+ _00113_ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12319__A1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11739__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ net257 _03950_ net1026 vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11790__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__B _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10291_ final_design.VGA_data_control.data_to_VGA\[23\] final_design.VGA_data_control.data_to_VGA\[22\]
+ final_design.VGA_data_control.data_to_VGA\[21\] final_design.VGA_data_control.data_to_VGA\[20\]
+ net1063 net1062 vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12030_ net1670 net226 net398 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold170 final_design.VGA_data_control.ready_data\[13\] vssd1 vssd1 vccd1 vccd1 net1523
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08113__S net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06422__A final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold181 final_design.cpu.reg_window\[718\] vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_151_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 final_design.cpu.reg_window\[252\] vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout650 _05946_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout661 net663 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_4
Xfanout672 _01503_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_4
Xfanout683 net684 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__buf_4
X_13981_ clknet_leaf_12_clk _01212_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[969\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout694 net695 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_4
XANTENNA__11474__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12932_ clknet_leaf_109_clk _00170_ net1214 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_166_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12867__Q final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12863_ clknet_leaf_82_clk _00101_ net1248 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14008__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11814_ net227 net1898 net268 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__mux2_1
XANTENNA__12255__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_164_Left_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ net218 net2193 net416 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12270__A3 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07399__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input95_X net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ net2528 net297 _06196_ net434 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_12_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13415_ clknet_leaf_6_clk _00646_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[403\]
+ sky130_fd_sc_hd__dfrtp_1
X_10627_ _05368_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13346_ clknet_leaf_21_clk _00577_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[334\]
+ sky130_fd_sc_hd__dfrtp_1
X_10558_ _05285_ _05303_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11781__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13277_ clknet_leaf_30_clk _00508_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[265\]
+ sky130_fd_sc_hd__dfrtp_1
X_10489_ net1054 final_design.reqhand.current_client\[1\] vssd1 vssd1 vccd1 vccd1
+ _05239_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_173_Left_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09726__A2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12228_ net580 _06156_ net511 net377 net1871 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12159_ net180 net2349 net387 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__mux2_1
XANTENNA__07832__S1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07862__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12089__A3 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11237__X _05941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11297__A1 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ final_design.cpu.reg_window\[472\] final_design.cpu.reg_window\[504\] net949
+ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__mux2_1
XANTENNA__12494__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06651_ final_design.cpu.reg_window\[346\] final_design.cpu.reg_window\[378\] net953
+ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09370_ _04286_ _04288_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__nand2_1
X_06582_ _01529_ _01530_ _01531_ _01532_ net788 net794 vssd1 vssd1 vccd1 vccd1 _01533_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_82_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08321_ final_design.cpu.reg_window\[136\] final_design.cpu.reg_window\[168\] net838
+ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12261__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06476__A1 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08252_ final_design.cpu.reg_window\[458\] final_design.cpu.reg_window\[490\] net854
+ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__mux2_1
XANTENNA__08870__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07203_ net769 _02153_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06957__A1_N net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08183_ _03132_ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__nor2_2
XFILLER_0_104_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07134_ final_design.cpu.reg_window\[715\] final_design.cpu.reg_window\[747\] net938
+ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__mux2_1
XANTENNA__10024__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07425__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06941__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08622__C1 _02156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07065_ final_design.cpu.reg_window\[525\] final_design.cpu.reg_window\[557\] net915
+ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__mux2_1
XANTENNA__07440__A3 _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout494_A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07772__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ final_design.cpu.reg_window\[977\] final_design.cpu.reg_window\[1009\] net836
+ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout759_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _03101_ _04497_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09272__B _04190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06918_ final_design.cpu.reg_window\[850\] final_design.cpu.reg_window\[882\] net904
+ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__mux2_1
XANTENNA__12485__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08689__C1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ _02845_ _02846_ _02847_ _02848_ net688 net709 vssd1 vssd1 vccd1 vccd1 _02849_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07587__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09350__B1 _04231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09637_ _04084_ _04264_ _04275_ _04073_ _04555_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a221o_1
X_06849_ final_design.cpu.reg_window\[148\] final_design.cpu.reg_window\[180\] net947
+ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1191_X net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout547_X net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07900__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12237__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ _04485_ _04486_ net476 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09102__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08519_ final_design.cpu.reg_window\[834\] final_design.cpu.reg_window\[866\] net866
+ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__mux2_1
XANTENNA__07113__C1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09499_ _02609_ _04050_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12252__A3 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06467__A1 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11323__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11530_ net1713 net186 net526 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__mux2_1
XANTENNA__06417__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09405__A1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11461_ net219 net2299 net307 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13200_ clknet_leaf_105_clk _00431_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[188\]
+ sky130_fd_sc_hd__dfrtp_1
X_10412_ _03321_ _05181_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__nor2_1
X_14180_ clknet_leaf_73_clk _01354_ net1246 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11392_ net740 _03811_ _06076_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11469__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13131_ clknet_leaf_13_clk _00362_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[119\]
+ sky130_fd_sc_hd__dfrtp_1
X_10343_ net1527 net1022 net999 final_design.data_from_mem\[28\] vssd1 vssd1 vccd1
+ vccd1 _00100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input55_A mem_adr_start[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ net2564 _05133_ net810 vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__o21ai_1
X_13062_ clknet_leaf_171_clk _00293_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08916__B1 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ _06215_ net292 net403 net2269 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__a22o_1
XANTENNA__11993__A _05869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09734__Y _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08401__A1_N net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10723__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout480 net482 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout491 net492 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11279__A1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10402__A _03481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12476__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13964_ clknet_leaf_122_clk _01195_ net1197 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[952\]
+ sky130_fd_sc_hd__dfrtp_1
X_12915_ clknet_leaf_33_clk _00153_ net1129 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
X_13895_ clknet_leaf_16_clk _01126_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[883\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09892__A1 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12228__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12846_ clknet_leaf_81_clk _00084_ net1247 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09644__A1 _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12243__A3 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11728_ net436 net590 _06222_ net297 net1545 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ net185 net641 vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12400__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold906 final_design.cpu.reg_window\[465\] vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold917 final_design.cpu.reg_window\[339\] vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 final_design.cpu.reg_window\[620\] vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ clknet_leaf_109_clk _00560_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[317\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09698__A2_N net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold939 final_design.cpu.reg_window\[385\] vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_36_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08870_ net632 _03817_ _03818_ net260 vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__a211o_1
XANTENNA__07805__S1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07821_ _02610_ _02642_ _02706_ _02771_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_32_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07591__C1 _02503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12467__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ net610 _02698_ _02674_ net559 vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__o211a_1
XANTENNA__10312__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07569__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06703_ final_design.cpu.reg_window\[537\] final_design.cpu.reg_window\[569\] net944
+ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__mux2_1
X_07683_ _02628_ _02633_ net720 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11842__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ net497 _04111_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__nand2_4
XANTENNA__12219__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11690__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06634_ final_design.cpu.reg_window\[795\] final_design.cpu.reg_window\[827\] net960
+ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__mux2_1
XANTENNA__06936__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09353_ net481 _04083_ _04086_ _04269_ _04271_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__o311a_1
XFILLER_0_19_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06565_ final_design.cpu.reg_window\[93\] final_design.cpu.reg_window\[125\] net959
+ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__mux2_1
XANTENNA__08438__A2 _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12234__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout242_A _05875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08304_ _03251_ _03252_ _03253_ _03254_ net688 net709 vssd1 vssd1 vccd1 vccd1 _03255_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06496_ final_design.cpu.reg_window\[670\] final_design.cpu.reg_window\[702\] net931
+ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__mux2_1
X_09284_ net614 _03549_ net562 _02422_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07110__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08235_ final_design.cpu.reg_window\[715\] final_design.cpu.reg_window\[747\] net856
+ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout507_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ net717 _03110_ net730 vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__o21a_1
XANTENNA__06671__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07117_ final_design.cpu.reg_window\[331\] final_design.cpu.reg_window\[363\] net938
+ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
XANTENNA__09267__B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08097_ final_design.cpu.reg_window\[12\] final_design.cpu.reg_window\[44\] net846
+ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1037_X net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07048_ final_design.data_from_mem\[14\] net982 _01997_ vssd1 vssd1 vccd1 vccd1 _01999_
+ sky130_fd_sc_hd__o21ai_4
Xclkload90 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout876_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08374__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08999_ _02452_ _02454_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10961_ net52 _05688_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net1064 _06340_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13680_ clknet_leaf_105_clk _00911_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[668\]
+ sky130_fd_sc_hd__dfrtp_1
X_10892_ _05600_ _05621_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__nor2_1
X_12631_ final_design.VGA_data_control.ready_data\[3\] net1032 net987 final_design.data_from_mem\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12225__A3 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08346__B net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12562_ _06225_ net349 net324 net2023 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11513_ net2143 net213 net526 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12493_ _06153_ net357 net333 net1674 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14232_ net1297 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_135_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11444_ net436 _06094_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11197__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12880__Q final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ clknet_leaf_82_clk net1717 net1242 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09177__B _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11375_ net670 _03826_ net748 vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13114_ clknet_leaf_164_clk _00345_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[102\]
+ sky130_fd_sc_hd__dfrtp_1
X_10326_ net1469 net1024 net1001 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1
+ vccd1 _00083_ sky130_fd_sc_hd__a22o_1
X_14094_ clknet_leaf_83_clk _01291_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13045_ clknet_leaf_40_clk _00276_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[33\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_2__f_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__09157__A3 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10257_ final_design.uart.BAUD_counter\[21\] _05123_ vssd1 vssd1 vccd1 vccd1 _05124_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09905__B _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1220 net1224 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_147_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09193__A _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1231 net1234 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__clkbuf_4
X_10188_ _05072_ _05077_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__or2_2
Xfanout1242 net1243 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_4
Xfanout1253 net1254 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09314__A0 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13947_ clknet_leaf_154_clk _01178_ net1118 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[935\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06679__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10475__A2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ clknet_leaf_126_clk _01109_ net1192 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[866\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06756__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12829_ net1369 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09078__C1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09617__A1 _04066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12216__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11975__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_150_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_150_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08020_ _02967_ _02968_ _02969_ _02970_ net683 net705 vssd1 vssd1 vccd1 vccd1 _02971_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold703 final_design.cpu.reg_window\[174\] vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 final_design.cpu.reg_window\[582\] vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold725 final_design.cpu.reg_window\[569\] vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold736 final_design.cpu.reg_window\[864\] vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold747 final_design.cpu.reg_window\[396\] vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 final_design.cpu.reg_window\[988\] vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07800__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold769 final_design.cpu.reg_window\[509\] vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ net265 _04889_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__nand2_1
XANTENNA__11837__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08922_ _02465_ _02466_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08853_ _03803_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout192_A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11138__A _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07804_ final_design.cpu.reg_window\[921\] final_design.cpu.reg_window\[953\] net860
+ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__mux2_1
X_08784_ final_design.CPU_instr_adr\[12\] _02064_ _03734_ vssd1 vssd1 vccd1 vccd1
+ _03735_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_169_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07735_ net723 _02679_ net731 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__o21a_1
XANTENNA__12668__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09856__A1 _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__A2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07666_ final_design.cpu.reg_window\[94\] final_design.cpu.reg_window\[126\] net847
+ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__mux2_1
XANTENNA__06666__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ net451 _04322_ _04323_ _04321_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_49_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06617_ final_design.reqhand.instruction\[28\] final_design.data_from_mem\[28\] net983
+ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__mux2_2
XFILLER_0_137_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12207__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07597_ final_design.cpu.reg_window\[413\] final_design.cpu.reg_window\[445\] net883
+ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09336_ _02673_ _03602_ _04254_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__or3_1
X_06548_ net751 net674 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11966__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09267_ net73 net74 _04185_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_141_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_141_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06479_ _01423_ _01424_ _01428_ _01429_ net779 net800 vssd1 vssd1 vccd1 vccd1 _01430_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1154_X net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09278__A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08218_ final_design.cpu.reg_window\[331\] final_design.cpu.reg_window\[363\] net857
+ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09198_ net497 _04054_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__nand2_2
XANTENNA__11179__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11718__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08149_ net620 _03096_ _03098_ net544 vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_30_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09792__A0 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11160_ final_design.data_from_mem\[2\] net253 _05855_ _05872_ vssd1 vssd1 vccd1
+ vccd1 _05873_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11747__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10111_ final_design.VGA_data_control.v_count\[2\] _05019_ final_design.VGA_data_control.v_count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_8_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11091_ _05799_ _05810_ _05812_ net59 vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09139__A3 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _04198_ _04253_ _04329_ _04960_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__and4_1
XANTENNA__06430__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 final_design.cpu.reg_window\[19\] vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 final_design.cpu.reg_window\[31\] vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 final_design.reqhand.instruction\[18\] vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 final_design.VGA_data_control.data_to_VGA\[2\] vssd1 vssd1 vccd1 vccd1 net1416
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold74 net152 vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 final_design.VGA_data_control.data_to_VGA\[20\] vssd1 vssd1 vccd1 vccd1 net1438
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 net107 vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ clknet_leaf_86_clk _01032_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[789\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10887__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ _05869_ net242 net636 vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__and3_1
XANTENNA__11482__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_10__f_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13732_ clknet_leaf_98_clk _00963_ net1227 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[720\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10944_ _05542_ _05603_ _05668_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__or3_1
XANTENNA__11654__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10457__A2 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08357__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12875__Q final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07261__A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13663_ clknet_leaf_133_clk _00894_ net1166 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[651\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10875_ _05602_ _05605_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12614_ net1398 final_design.reqhand.data_from_UART\[0\] _05080_ vssd1 vssd1 vccd1
+ vccd1 _01307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13594_ clknet_leaf_160_clk _00825_ net1105 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[582\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12545_ _06208_ net351 net324 net2105 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_132_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_152_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08804__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06833__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09188__A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12476_ _06136_ net353 net333 net2195 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07200__S net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ net1284 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_124_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11427_ net2032 net203 net311 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__mux2_1
XANTENNA_5 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09475__X _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ clknet_leaf_77_clk _01320_ net1255 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ net668 _03840_ net740 vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10393__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10309_ net1061 _05155_ _05157_ _05162_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__o31ai_1
X_14077_ clknet_leaf_43_clk _01274_ net1153 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10414__X _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11289_ _01909_ net649 _05985_ _05986_ net662 vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_5_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13028_ clknet_leaf_93_clk _00259_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11342__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1050 _01410_ vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_4
Xfanout1061 final_design.VGA_data_control.h_count\[4\] vssd1 vssd1 vccd1 vccd1 net1061
+ sky130_fd_sc_hd__buf_2
Xfanout1072 final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1 net1072
+ sky130_fd_sc_hd__clkbuf_4
Xfanout1083 net1104 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_4
Xfanout1094 net1095 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__buf_2
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09838__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07520_ _01662_ _02470_ _01631_ _01632_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07451_ final_design.cpu.reg_window\[0\] final_design.cpu.reg_window\[32\] net944
+ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07382_ final_design.cpu.reg_window\[322\] final_design.cpu.reg_window\[354\] net947
+ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09121_ net1006 net1004 vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__nor2_2
XANTENNA__07077__A1 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11948__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_123_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_44_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09052_ final_design.CPU_instr_adr\[9\] _03787_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_96_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06515__A final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08206__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08003_ _02950_ _02951_ _02952_ _02953_ net696 net715 vssd1 vssd1 vccd1 vccd1 _02954_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold500 final_design.cpu.reg_window\[560\] vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold511 final_design.cpu.reg_window\[362\] vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 final_design.cpu.reg_window\[966\] vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold533 final_design.cpu.reg_window\[577\] vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09826__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold544 final_design.cpu.reg_window\[995\] vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06588__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold555 final_design.cpu.reg_window\[565\] vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 final_design.cpu.reg_window\[775\] vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11581__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07785__C1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold577 final_design.cpu.reg_window\[266\] vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 final_design.cpu.reg_window\[642\] vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09954_ _03486_ net441 _04872_ net451 vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a211o_1
XANTENNA__11794__C net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold599 final_design.cpu.reg_window\[387\] vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1114_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08905_ net633 _03847_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__nor2_1
X_09885_ _03522_ _03640_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__xor2_1
Xhold1200 _00030_ vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout574_A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1211 final_design.uart.BAUD_counter\[27\] vssd1 vssd1 vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout195_X net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1222 final_design.reqhand.instruction\[4\] vssd1 vssd1 vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ final_design.CPU_instr_adr\[8\] _03786_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08767_ final_design.CPU_instr_adr\[0\] _02425_ _03716_ _03714_ vssd1 vssd1 vccd1
+ vccd1 _03718_ sky130_fd_sc_hd__a31o_1
XANTENNA__09829__A1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07718_ _01599_ net611 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__and2_1
XANTENNA__11636__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_68_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08698_ _01486_ _03646_ _03648_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_68_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07081__A _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07935__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07649_ _02596_ _02597_ _02598_ _02599_ net694 net702 vssd1 vssd1 vccd1 vccd1 _02600_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ _05400_ _05401_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__nand2_1
XANTENNA__08905__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11939__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09319_ net532 net455 vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10591_ _05315_ _05318_ _05335_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_114_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12330_ net680 net658 _06268_ net363 net1608 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__a32o_1
XFILLER_0_106_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06910__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ net581 _06190_ net512 net373 net1431 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08112__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14000_ clknet_leaf_112_clk _01231_ net1211 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[988\]
+ sky130_fd_sc_hd__dfrtp_1
X_11212_ net652 _05918_ _05916_ net663 vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a211o_1
XANTENNA__07955__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12192_ net1972 net183 net383 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__mux2_1
XANTENNA__10375__B2 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ _04939_ net660 net600 _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__o211a_1
X_11074_ _05793_ _05794_ _05796_ net1046 net1382 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__a32o_1
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10025_ _04108_ _04398_ net319 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12419__A3 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12101__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ _06178_ net278 net404 net1883 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__a22o_1
XANTENNA__10410__A _03352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13715_ clknet_leaf_35_clk _00946_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[703\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ _05654_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13646_ clknet_leaf_117_clk _00877_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[634\]
+ sky130_fd_sc_hd__dfrtp_1
X_10858_ _05588_ _05589_ _05568_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_144_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12052__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13577_ clknet_leaf_85_clk _00808_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[565\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_105_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10789_ _05508_ _05524_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08351__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10602__A2 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12528_ _06190_ net350 net328 net1678 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ net1700 net185 net338 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12355__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10366__B2 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06989__B _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14129_ clknet_leaf_74_clk final_design.vga.v_next_state\[0\] net1245 vssd1 vssd1
+ vccd1 vccd1 final_design.vga.v_current_state\[0\] sky130_fd_sc_hd__dfrtp_1
Xfanout309 net310 vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_8
XANTENNA__07782__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13172__CLK clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06951_ final_design.cpu.reg_window\[721\] final_design.cpu.reg_window\[753\] net910
+ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__mux2_1
XANTENNA__11315__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09652__Y _04571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _02804_ net446 net443 _02800_ _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__o221a_1
XANTENNA__11866__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06882_ final_design.cpu.reg_window\[19\] final_design.cpu.reg_window\[51\] net908
+ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08621_ _03198_ _03571_ _03570_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__a21oi_1
X_08552_ final_design.cpu.reg_window\[961\] final_design.cpu.reg_window\[993\] net851
+ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__mux2_1
XANTENNA__11618__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07503_ _01969_ _01970_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_46_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08483_ final_design.cpu.reg_window\[195\] final_design.cpu.reg_window\[227\] net861
+ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__mux2_1
XANTENNA__12291__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07434_ final_design.cpu.reg_window\[577\] final_design.cpu.reg_window\[609\] net932
+ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__mux2_1
XANTENNA__08590__S0 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12973__RESET_B net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07365_ final_design.cpu.reg_window\[899\] final_design.cpu.reg_window\[931\] net942
+ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout322_A _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09104_ _02430_ _04024_ _04025_ net628 vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11151__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09259__C net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07296_ _02243_ _02244_ _02245_ _02246_ net774 net795 vssd1 vssd1 vccd1 vccd1 _02247_
+ sky130_fd_sc_hd__mux4_1
X_09035_ _03963_ _03965_ net258 vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1231_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout208_X net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07775__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12346__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold330 final_design.cpu.reg_window\[834\] vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 final_design.cpu.reg_window\[733\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10357__B2 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold352 final_design.cpu.reg_window\[562\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout691_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold363 final_design.VGA_data_control.data_to_VGA\[22\] vssd1 vssd1 vccd1 vccd1 net1716
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09275__B net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 final_design.cpu.reg_window\[60\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 final_design.cpu.reg_window\[903\] vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 final_design.cpu.reg_window\[753\] vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 net812 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__buf_2
Xfanout821 net823 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_4
Xfanout832 net834 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_4
X_09937_ _03388_ net439 _04109_ _04309_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__o221a_1
Xfanout843 net845 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_4
Xfanout854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__buf_4
XANTENNA_fanout956_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout865 net867 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout876 net877 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__buf_2
Xfanout887 _01818_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_4
X_09868_ net737 _04772_ _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__and3_1
Xhold1030 final_design.cpu.reg_window\[103\] vssd1 vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11857__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout898 net899 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__clkbuf_8
Xhold1041 final_design.cpu.reg_window\[110\] vssd1 vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ _03668_ _03769_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__nor2_1
Xhold1052 final_design.cpu.reg_window\[635\] vssd1 vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 final_design.cpu.reg_window\[948\] vssd1 vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 final_design.cpu.reg_window\[115\] vssd1 vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ _03455_ _03557_ _03560_ _03457_ _03424_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__o311a_1
XANTENNA__13008__RESET_B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08178__Y _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1085 final_design.cpu.reg_window\[124\] vssd1 vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ net200 net2270 net266 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__mux2_1
Xhold1096 final_design.cpu.reg_window\[627\] vssd1 vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_77_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07289__A1 _01628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ net188 net1902 net418 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__mux2_1
XANTENNA__11760__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13500_ clknet_leaf_147_clk _00731_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[488\]
+ sky130_fd_sc_hd__dfrtp_1
X_10712_ _05449_ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06854__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06707__X _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11692_ net582 net422 _06204_ net296 net1666 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_4_3__f_clk_X clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13431_ clknet_leaf_145_clk _00662_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[419\]
+ sky130_fd_sc_hd__dfrtp_1
X_10643_ _05362_ _05383_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10045__B1 _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input85_A memory_size[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13362_ clknet_leaf_27_clk _00593_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[350\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_172_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10574_ final_design.CPU_instr_adr\[6\] _05319_ net1067 vssd1 vssd1 vccd1 vccd1 _05320_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09450__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10596__B2 _01371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11793__B1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12313_ net1903 net221 net366 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_86_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13293_ clknet_leaf_141_clk _00524_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[281\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12337__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12244_ net578 _06174_ net500 net373 net1534 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__a32o_1
XANTENNA__11545__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12175_ net2486 net213 net382 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08961__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ _01487_ net665 net1030 vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_43_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10899__X _05629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11057_ net89 net1058 vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__nor2_1
XANTENNA__09913__B _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13431__RESET_B net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09910__B1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ _03642_ _04045_ _04089_ _03641_ _04926_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_95_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11236__A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07978__A1_N net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11959_ _06160_ net286 net405 net1948 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06617__X _01568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09140__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08229__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13629_ clknet_leaf_32_clk _00860_ net1129 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[617\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07150_ net542 _02098_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09928__X _04847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07081_ _02026_ _02031_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09729__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09376__A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10339__B2 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07204__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09744__A3 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_wire545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_14__f_clk_X clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07983_ net617 _02929_ _02931_ _01908_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a211o_1
XANTENNA__11845__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ net546 net545 net544 net543 net453 net462 vssd1 vssd1 vccd1 vccd1 _04641_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06934_ final_design.cpu.reg_window\[465\] final_design.cpu.reg_window\[497\] net918
+ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__mux2_1
XANTENNA__13172__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ net78 _04188_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06865_ _01381_ net1051 net1008 net1005 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout272_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ _03520_ _03521_ _03554_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_171_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09584_ _04144_ _04153_ _04154_ _04155_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_26_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06796_ final_design.cpu.reg_window\[918\] final_design.cpu.reg_window\[950\] net905
+ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08535_ net624 _03481_ _03482_ net532 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_49_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1181_A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout537_A _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07366__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08466_ _02297_ net625 vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_102_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12973__Q final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07417_ final_design.cpu.reg_window\[385\] final_design.cpu.reg_window\[417\] net930
+ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08397_ final_design.cpu.reg_window\[582\] final_design.cpu.reg_window\[614\] net830
+ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout704_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1067_X net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire529 _02731_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_4
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ _02294_ _02297_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10578__A1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07279_ final_design.cpu.reg_window\[966\] final_design.cpu.reg_window\[998\] net913
+ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1234_X net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09018_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__inv_2
X_10290_ final_design.VGA_data_control.data_to_VGA\[19\] final_design.VGA_data_control.data_to_VGA\[18\]
+ final_design.VGA_data_control.data_to_VGA\[17\] final_design.VGA_data_control.data_to_VGA\[16\]
+ net1063 net1062 vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__mux4_1
XANTENNA__08190__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09717__C _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13942__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold160 _01311_ vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 final_design.VGA_data_control.ready_data\[2\] vssd1 vssd1 vccd1 vccd1 net1524
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold182 final_design.cpu.reg_window\[94\] vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 final_design.cpu.reg_window\[219\] vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 net641 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_109_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout651 net653 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11755__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout662 net663 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_2
X_13980_ clknet_leaf_153_clk _01211_ net1118 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[968\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout673 net675 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_4
XANTENNA__06849__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout684 net698 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_4
Xfanout695 net698 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_4
X_12931_ clknet_leaf_110_clk _00169_ net1214 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11056__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12862_ clknet_leaf_82_clk _00100_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11813_ net242 net2286 net268 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12255__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08554__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ net220 net2346 net417 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12883__Q final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11675_ net588 net241 net636 vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ clknet_leaf_0_clk _00645_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[402\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12558__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10626_ net99 final_design.VGA_adr\[7\] vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__nand2_1
XANTENNA_input88_X net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11766__A0 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13345_ clknet_leaf_152_clk _00576_ net1116 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[333\]
+ sky130_fd_sc_hd__dfrtp_1
X_10557_ _05267_ _05285_ _05303_ _05283_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__o211a_1
XANTENNA__09908__B _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13276_ clknet_leaf_147_clk _00507_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[264\]
+ sky130_fd_sc_hd__dfrtp_1
X_10488_ net1031 net1073 vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09187__A1 _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12227_ net581 _06155_ net512 net377 net1760 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__a32o_1
XANTENNA__09726__A3 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09924__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ net183 net2278 net386 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__mux2_1
XANTENNA__06945__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ net1650 net1046 net1016 _05829_ vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12089_ net592 _06061_ net518 net395 net2244 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_34_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07444__A _02390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06650_ net560 _01599_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06581_ final_design.cpu.reg_window\[541\] final_design.cpu.reg_window\[573\] net957
+ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08320_ final_design.cpu.reg_window\[200\] final_design.cpu.reg_window\[232\] net838
+ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08251_ final_design.cpu.reg_window\[266\] final_design.cpu.reg_window\[298\] net854
+ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07202_ _02149_ _02150_ _02151_ _02152_ net780 net799 vssd1 vssd1 vccd1 vccd1 _02153_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12549__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14255__1320 vssd1 vssd1 vccd1 vccd1 _14255__1320/HI net1320 sky130_fd_sc_hd__conb_1
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08182_ net616 _03129_ _03131_ _01966_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_132_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11757__A0 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07133_ _02080_ _02081_ _02082_ _02083_ net783 net802 vssd1 vssd1 vccd1 vccd1 _02084_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07425__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08722__B _01881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07064_ final_design.cpu.reg_window\[589\] final_design.cpu.reg_window\[621\] net915
+ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1027_A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout487_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06669__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ net725 _02916_ net730 vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09045__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ _03102_ net446 _04617_ _04623_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__o211a_1
X_06917_ net767 _01867_ net754 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07036__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08689__B1 _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07897_ final_design.cpu.reg_window\[151\] final_design.cpu.reg_window\[183\] net843
+ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout654_A _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09350__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ _04107_ _04277_ _04116_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_104_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07587__S1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06848_ final_design.cpu.reg_window\[212\] final_design.cpu.reg_window\[244\] net949
+ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07361__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ net554 net553 net552 net551 net453 net462 vssd1 vssd1 vccd1 vccd1 _04486_
+ sky130_fd_sc_hd__mux4_1
X_06779_ _01726_ _01727_ _01728_ _01729_ net774 net795 vssd1 vssd1 vccd1 vccd1 _01730_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout919_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ net721 _03462_ net731 vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__o21a_1
XANTENNA__11604__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09498_ _04074_ _04403_ _04416_ _04400_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__o211a_1
XFILLER_0_136_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11996__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08310__C1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08449_ final_design.cpu.reg_window\[132\] final_design.cpu.reg_window\[164\] net858
+ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__mux2_1
XANTENNA__11323__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ net219 net646 vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11748__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_clk_X clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10411_ net255 _05188_ net1040 net1618 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11212__A2 _05918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11391_ net668 _03807_ net740 vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13130_ clknet_leaf_0_clk _00361_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10420__B1 _05193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10342_ net1509 net1024 net1001 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1
+ vccd1 _00099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08124__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13061_ clknet_leaf_4_clk _00292_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_10273_ final_design.uart.BAUD_counter\[27\] _05133_ vssd1 vssd1 vccd1 vccd1 _05134_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08916__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07719__A2 _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ _06214_ net290 net402 net2189 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__a22o_1
XANTENNA__11993__B net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_A mem_adr_start[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11920__A0 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10723__B2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout470 _03518_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_2
Xfanout481 net482 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_2
XANTENNA__12878__Q final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout492 net495 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_2
X_13963_ clknet_leaf_15_clk _01194_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[951\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10402__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_85_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12914_ clknet_leaf_156_clk _00152_ net1114 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
X_13894_ clknet_leaf_165_clk _01125_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[882\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12845_ clknet_leaf_80_clk _00083_ net1249 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12228__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06608__A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11987__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11727_ net182 net636 vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11658_ net589 net423 _06186_ net301 net1465 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11739__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10609_ _05351_ _05352_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__nor2_1
XANTENNA__07407__A1 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09638__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11589_ net591 net423 _06150_ net305 net1707 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__a32o_1
XFILLER_0_12_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold907 final_design.cpu.reg_window\[527\] vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold918 final_design.cpu.reg_window\[433\] vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ clknet_leaf_113_clk _00559_ net1212 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[316\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10411__B1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold929 final_design.cpu.reg_window\[422\] vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13259_ clknet_leaf_15_clk _00490_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[247\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07873__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11248__X _05951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ _02734_ _02736_ _02766_ _02767_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__o22a_1
XANTENNA__09373__B _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07174__A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ net559 _02700_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__or2_2
XFILLER_0_159_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12467__A1 _06127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_76_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06702_ final_design.cpu.reg_window\[601\] final_design.cpu.reg_window\[633\] net940
+ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__mux2_1
XANTENNA__07569__S1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09660__Y _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07682_ _02629_ _02630_ _02631_ _02632_ net687 net701 vssd1 vssd1 vccd1 vccd1 _02633_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09421_ net498 _04112_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__nor2_1
X_06633_ final_design.cpu.reg_window\[859\] final_design.cpu.reg_window\[891\] net960
+ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09352_ _02673_ net447 net444 _02670_ _04270_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__o221a_1
XANTENNA__09096__B1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06564_ _01511_ _01512_ _01513_ _01514_ net788 net806 vssd1 vssd1 vccd1 vccd1 _01515_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08677__A_N net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11978__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08303_ final_design.cpu.reg_window\[905\] final_design.cpu.reg_window\[937\] net842
+ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_150_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09283_ _04200_ _04201_ net476 vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__mux2_1
X_06495_ final_design.cpu.reg_window\[734\] final_design.cpu.reg_window\[766\] net931
+ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ _03181_ _03182_ _03183_ _03184_ net691 net711 vssd1 vssd1 vccd1 vccd1 _03185_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06952__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08165_ net725 _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout402_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1144_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07116_ _02065_ _02066_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_165_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08096_ final_design.cpu.reg_window\[76\] final_design.cpu.reg_window\[108\] net846
+ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload80 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__clkinv_4
X_07047_ final_design.data_from_mem\[14\] net982 _01997_ vssd1 vssd1 vccd1 vccd1 _01998_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload91 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__inv_6
XFILLER_0_140_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12155__A0 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11902__A0 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout771_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__A2 _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10503__A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ net630 _03932_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__nor2_1
X_07949_ _02897_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__or2_2
XFILLER_0_173_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_67_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ net678 _05674_ _05687_ net978 _05686_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__o221a_1
XFILLER_0_173_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09619_ _04077_ net320 vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__nand2_1
X_10891_ _05621_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12630_ _06302_ net1416 net992 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__mux2_1
XANTENNA__09087__A0 final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11969__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12561_ _06224_ net350 net324 net1710 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07958__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11512_ net1847 net216 net525 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__mux2_1
XANTENNA__09739__A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12492_ _06152_ _06277_ net334 net2136 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14231_ net1296 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11443_ net681 net648 vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__and2_2
XFILLER_0_117_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09458__B net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11197__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14162_ clknet_leaf_82_clk _01336_ net1243 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11374_ net438 net596 _06061_ net318 net1658 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_169_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13113_ clknet_leaf_167_clk _00344_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[101\]
+ sky130_fd_sc_hd__dfrtp_1
X_10325_ net1543 net1024 net1001 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1
+ vccd1 _00082_ sky130_fd_sc_hd__a22o_1
X_14093_ clknet_leaf_82_clk _01290_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_13044_ clknet_leaf_102_clk _00275_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_10256_ _05123_ net810 _05122_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__and3b_1
Xfanout1210 net1216 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__clkbuf_4
Xfanout1221 net1222 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09193__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1232 net1234 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12104__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ _05073_ _05074_ _05075_ _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__or4_1
Xfanout1243 net1256 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__buf_2
Xfanout1254 net1255 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12449__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09314__A1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08117__A2 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13946_ clknet_leaf_163_clk _01177_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[934\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13877_ clknet_leaf_24_clk _01108_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[865\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11244__A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ net1359 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12621__A1 final_design.reqhand.data_from_UART\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12759_ net967 _06382_ _06394_ _06395_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07868__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold704 final_design.cpu.reg_window\[246\] vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold715 final_design.cpu.reg_window\[930\] vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 final_design.cpu.reg_window\[192\] vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold737 final_design.cpu.reg_window\[334\] vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold748 final_design.cpu.reg_window\[793\] vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07800__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09970_ _03327_ net447 _04119_ _04066_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__o221a_1
Xhold759 final_design.cpu.reg_window\[391\] vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08921_ _03757_ _03863_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__xor2_1
XANTENNA__12998__RESET_B net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08852_ final_design.CPU_instr_adr\[31\] _03802_ vssd1 vssd1 vccd1 vccd1 _03803_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_51_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07175__Y _02126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11360__A1 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ final_design.cpu.reg_window\[985\] final_design.cpu.reg_window\[1017\] net859
+ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08783_ _03688_ _03732_ _03687_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__and3b_1
Xclkbuf_leaf_49_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout185_A _06060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07734_ net728 _02684_ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_140_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06947__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07632__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07665_ _02612_ _02613_ _02614_ _02615_ net689 net708 vssd1 vssd1 vccd1 vccd1 _02616_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout352_A _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ _02606_ _04171_ _02576_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1094_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06616_ net898 _01559_ _01565_ _01547_ _01553_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__a32o_4
XANTENNA__09069__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07596_ final_design.cpu.reg_window\[477\] final_design.cpu.reg_window\[509\] net883
+ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ _02704_ _04049_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06547_ _01484_ _01488_ net746 _01494_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__or4_1
XANTENNA__10993__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12684__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12612__B2 final_design.data_from_mem\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_X net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09266_ net72 _04184_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__or2_2
XFILLER_0_118_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06682__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06478_ final_design.cpu.reg_window\[414\] final_design.cpu.reg_window\[446\] net930
+ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08217_ _02097_ net615 vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09197_ net499 _04055_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__nor2_2
XFILLER_0_31_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08148_ net604 _03096_ _03072_ _02026_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__o211a_1
XANTENNA__08044__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09792__A1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08079_ _02994_ _02995_ _03025_ _03027_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_112_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10110_ final_design.VGA_data_control.v_count\[2\] final_design.VGA_data_control.v_count\[3\]
+ _05019_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_8_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11090_ net975 _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12679__B2 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06711__A _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ _04479_ _04532_ _04552_ _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__and4_1
XANTENNA__11351__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 final_design.cpu.reg_window\[17\] vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 final_design.reqhand.instruction\[16\] vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 final_design.reqhand.instruction\[23\] vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 final_design.uart.working_data\[2\] vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 final_design.reqhand.instruction\[11\] vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11763__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold75 net157 vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 final_design.reqhand.instruction\[28\] vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ clknet_leaf_119_clk _01031_ net1199 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[788\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold97 final_design.VGA_data_control.data_to_VGA\[15\] vssd1 vssd1 vccd1 vccd1 net1450
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ _06195_ net286 net401 net1969 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__a22o_1
X_10943_ _05604_ _05668_ _05669_ _05670_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__o211ai_1
X_13731_ clknet_leaf_2_clk _00962_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[719\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11654__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07261__B _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10874_ _05602_ _05605_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__or2_1
Xclkbuf_3_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_clk sky130_fd_sc_hd__clkbuf_8
X_13662_ clknet_leaf_149_clk _00893_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[650\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12613_ net1995 net1009 net995 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1
+ vccd1 _01306_ sky130_fd_sc_hd__a22o_1
X_13593_ clknet_leaf_167_clk _00824_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[581\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12603__B2 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09469__A _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10614__B1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12544_ _06207_ net347 net324 net1668 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06592__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12891__Q final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12475_ _06135_ net348 net331 net2073 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__a22o_1
XANTENNA__10408__A _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14214_ net1283 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XFILLER_0_22_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11426_ net1633 net222 net314 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14145_ clknet_leaf_77_clk _01319_ net1254 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11357_ net591 net423 _06046_ net317 net2315 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09916__B _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10393__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ _05147_ _05159_ _05161_ final_design.VGA_data_control.h_count\[5\] vssd1
+ vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14076_ clknet_leaf_52_clk _01273_ net1153 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11288_ net743 _03918_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__nand2_1
X_13027_ clknet_leaf_7_clk _00258_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08338__A2 _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10239_ final_design.uart.BAUD_counter\[13\] final_design.uart.BAUD_counter\[14\]
+ _05109_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__and3_1
XANTENNA__11342__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1040 net1044 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__buf_4
Xfanout1051 _01394_ vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_2
Xfanout1062 final_design.VGA_data_control.h_count\[2\] vssd1 vssd1 vccd1 vccd1 net1062
+ sky130_fd_sc_hd__clkbuf_4
Xfanout1073 final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1 net1073
+ sky130_fd_sc_hd__buf_2
Xfanout1084 net1085 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__clkbuf_4
Xfanout1095 net1104 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08548__A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13929_ clknet_leaf_86_clk _01160_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[917\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10853__A0 final_design.CPU_instr_adr\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07450_ final_design.cpu.reg_window\[64\] final_design.cpu.reg_window\[96\] net944
+ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06521__A1 final_design.data_from_mem\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07381_ _02325_ _02330_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09120_ net975 _04037_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07598__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12070__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09051_ net631 _03979_ _03977_ net258 vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08002_ final_design.cpu.reg_window\[912\] final_design.cpu.reg_window\[944\] net878
+ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__mux2_1
XANTENNA__12358__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold501 final_design.cpu.reg_window\[378\] vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10908__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10908__B2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold512 final_design.cpu.reg_window\[559\] vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 final_design.cpu.reg_window\[781\] vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 final_design.cpu.reg_window\[589\] vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09826__B _04744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold545 final_design.cpu.reg_window\[323\] vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06588__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06802__Y _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold556 final_design.cpu.reg_window\[545\] vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08730__B _02000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11581__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 final_design.cpu.reg_window\[886\] vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 final_design.cpu.reg_window\[905\] vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 final_design.cpu.reg_window\[70\] vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _03487_ net444 vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_115_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09526__A1 _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11149__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08904_ _01661_ _01662_ _02469_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__o21ai_1
X_09884_ _04789_ _04791_ _04792_ _04802_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__and4bb_1
XANTENNA_fanout1107_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1201 net115 vssd1 vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11333__B2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1212 final_design.CPU_instr_adr\[13\] vssd1 vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ final_design.CPU_instr_adr\[7\] final_design.CPU_instr_adr\[6\] _03785_ vssd1
+ vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__and3_1
XANTENNA__10988__A _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout567_A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout188_X net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ _03714_ _03716_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__and2b_1
XANTENNA__06677__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09829__A2 _04744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07717_ net893 _02649_ _02655_ _02661_ _02667_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__o32a_4
XANTENNA__13967__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11155__Y _05869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08697_ _02028_ _02062_ _01998_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout734_A _01493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07935__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07648_ final_design.cpu.reg_window\[540\] final_design.cpu.reg_window\[572\] net871
+ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ final_design.cpu.reg_window\[735\] final_design.cpu.reg_window\[767\] net846
+ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__mux2_1
XANTENNA__08464__Y _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09318_ net531 net459 vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_157_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10590_ _05311_ _05333_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09249_ _02735_ _02768_ _02766_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12349__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12260_ net592 _06189_ net518 net375 net1694 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ final_design.data_from_mem\[8\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__11758__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08112__S1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08568__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ net2076 net184 net383 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11142_ _05855_ _05856_ _05852_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a21o_1
XANTENNA__07537__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07871__S0 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11073_ net1018 _05795_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12521__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _02835_ net443 net440 _02834_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__o22a_1
XANTENNA__09752__A _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__Q final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11975_ _06177_ net280 net404 net2259 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__a22o_1
XANTENNA__10410__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13714_ clknet_leaf_41_clk _00945_ net1150 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[702\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10926_ _05632_ _05634_ _05652_ _05653_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10857_ net80 net1056 vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__nor2_1
X_13645_ clknet_leaf_137_clk _00876_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[633\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_160_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10788_ _05522_ _05523_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ clknet_leaf_126_clk _00807_ net1192 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[564\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10451__A1_N net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08351__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12527_ _06189_ net358 net330 net1993 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08831__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12458_ net2203 net187 net337 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11409_ net681 net438 _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12389_ net2005 net189 net272 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__mux2_1
XANTENNA__11563__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14128_ clknet_leaf_76_clk final_design.vga.v_next_count\[8\] net1252 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_123_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06950_ _01897_ _01898_ _01899_ _01900_ net778 net798 vssd1 vssd1 vccd1 vccd1 _01901_
+ sky130_fd_sc_hd__mux4_1
X_14059_ clknet_leaf_47_clk _00021_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12512__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06881_ final_design.cpu.reg_window\[83\] final_design.cpu.reg_window\[115\] net908
+ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__mux2_1
XANTENNA__11866__A2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08620_ _02127_ _03226_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__and2_1
X_08551_ final_design.cpu.reg_window\[769\] final_design.cpu.reg_window\[801\] net849
+ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__mux2_1
XANTENNA__11618__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07502_ _01970_ _02001_ _01969_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13378__RESET_B net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08482_ final_design.cpu.reg_window\[3\] final_design.cpu.reg_window\[35\] net864
+ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07433_ final_design.cpu.reg_window\[641\] final_design.cpu.reg_window\[673\] net936
+ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08590__S1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07364_ final_design.cpu.reg_window\[963\] final_design.cpu.reg_window\[995\] net942
+ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09103_ _03713_ _03718_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__xor2_1
XANTENNA__10054__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07295_ final_design.cpu.reg_window\[133\] final_design.cpu.reg_window\[165\] net904
+ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout315_A _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09034_ _03789_ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12942__RESET_B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 final_design.cpu.reg_window\[898\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold331 final_design.cpu.reg_window\[927\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12263__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1224_A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 final_design.cpu.reg_window\[698\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 final_design.cpu.reg_window\[550\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold364 _01337_ vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 final_design.uart.BAUD_counter\[22\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout800 net801 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_4
Xhold386 final_design.cpu.reg_window\[774\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout811 net812 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold397 final_design.cpu.reg_window\[61\] vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08970__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout822 net823 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_4
X_09936_ _03391_ net447 net444 _03389_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__o22a_1
Xfanout833 net834 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_2
Xfanout844 net845 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_4
Xfanout855 net887 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__buf_4
XANTENNA__12503__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07791__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout866 net867 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07605__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout851_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11857__A2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout877 net887 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__buf_2
X_09867_ _04125_ _04785_ _04784_ _04777_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a211o_1
Xhold1020 final_design.cpu.reg_window\[335\] vssd1 vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 net890 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__buf_8
XANTENNA_fanout949_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1031 final_design.cpu.reg_window\[889\] vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 net900 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11607__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1042 final_design.cpu.reg_window\[1014\] vssd1 vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ final_design.CPU_instr_adr\[24\] _01691_ vssd1 vssd1 vccd1 vccd1 _03769_
+ sky130_fd_sc_hd__nor2_1
Xhold1053 final_design.cpu.reg_window\[566\] vssd1 vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10511__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1064 final_design.cpu.reg_window\[514\] vssd1 vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ _04072_ _04714_ _04716_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__or3b_1
Xhold1075 final_design.cpu.reg_window\[430\] vssd1 vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 final_design.cpu.reg_window\[609\] vssd1 vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1097 final_design.cpu.reg_window\[369\] vssd1 vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08749_ final_design.CPU_instr_adr\[6\] _02240_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ net191 net2230 net418 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09683__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10711_ _05425_ _05429_ _05427_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11691_ net216 net635 vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10642_ _05364_ _05383_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__and2_2
XFILLER_0_153_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13430_ clknet_leaf_129_clk _00661_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[418\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13361_ clknet_leaf_111_clk _00592_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[349\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10573_ _05317_ _05318_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10596__A2 _05239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ net2223 net206 net364 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13292_ clknet_leaf_121_clk _00523_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[280\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input78_A memory_size[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08651__A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09738__A1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12243_ net574 _06173_ net509 net372 net1549 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11545__A1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ net1785 net215 net380 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__mux2_1
XANTENNA__07844__S0 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11125_ net816 _05839_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__and2_2
X_11056_ net88 net1058 net89 vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__or3b_1
XANTENNA__11848__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09910__A1 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10007_ _03640_ net440 vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__nor2_1
XANTENNA__10421__A _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12112__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11236__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11958_ net2144 net406 _06256_ net230 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__a22o_1
XANTENNA__09674__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06488__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ final_design.CPU_instr_adr\[22\] net1013 vssd1 vssd1 vccd1 vccd1 _05639_
+ sky130_fd_sc_hd__nor2_1
X_11889_ net240 net2297 net276 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08229__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13628_ clknet_leaf_152_clk _00859_ net1117 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[616\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09426__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13559_ clknet_leaf_144_clk _00790_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[547\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07876__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09657__A _04190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07080_ _02030_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08561__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09944__X _04863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07982_ net617 _02929_ _02931_ _01908_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__a211oi_2
X_06933_ _01883_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__inv_2
X_09721_ _03069_ net442 vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09652_ net449 _04569_ _04566_ net737 vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__o211ai_4
X_06864_ net898 _01796_ _01802_ _01808_ _01814_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__o32a_4
XANTENNA__08260__S0 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08603_ net614 _03550_ _03524_ _02419_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__o211ai_4
X_09583_ net322 _04500_ _04501_ _04494_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_171_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06795_ final_design.cpu.reg_window\[982\] final_design.cpu.reg_window\[1014\] net905
+ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08534_ net622 _03481_ _03482_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08465_ _02297_ net612 vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_102_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout432_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1174_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07140__B2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07416_ final_design.cpu.reg_window\[449\] final_design.cpu.reg_window\[481\] net930
+ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09417__A0 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12016__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ final_design.cpu.reg_window\[646\] final_design.cpu.reg_window\[678\] net830
+ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07347_ _02294_ _02297_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11224__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07278_ final_design.cpu.reg_window\[774\] final_design.cpu.reg_window\[806\] net917
+ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__mux2_1
XANTENNA__06690__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09017_ _03790_ _03949_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout899_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold150 final_design.cpu.reg_window\[710\] vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09854__X _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 final_design.VGA_data_control.ready_data\[21\] vssd1 vssd1 vccd1 vccd1 net1514
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 final_design.VGA_data_control.ready_data\[19\] vssd1 vssd1 vccd1 vccd1 net1525
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold183 final_design.cpu.reg_window\[187\] vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 final_design.VGA_data_control.data_to_VGA\[4\] vssd1 vssd1 vccd1 vccd1 net1547
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout630 _02506_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__buf_2
Xfanout641 _06157_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout652 net653 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_2
X_09919_ net488 _04646_ _04224_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_109_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout663 _05142_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08410__S net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout674 net675 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__buf_2
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout685 net686 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_3_1_0_clk_X clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12930_ clknet_leaf_90_clk _00168_ net1232 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dfrtp_1
Xfanout696 net697 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__buf_4
XANTENNA__11160__C1 _05872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06706__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07026__S net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ clknet_leaf_79_clk _00099_ net1249 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11812_ net228 net2070 net267 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__mux2_1
XANTENNA__08003__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07550__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08554__S1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11743_ net245 net2186 net417 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12007__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11674_ net430 net581 _06195_ net296 net2010 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_12_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ clknet_leaf_18_clk _00644_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[401\]
+ sky130_fd_sc_hd__dfrtp_1
X_10625_ net99 final_design.VGA_adr\[7\] vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14088__RESET_B net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10556_ net63 _05301_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__xnor2_1
X_13344_ clknet_leaf_39_clk _00575_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[332\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ _05235_ _05236_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__nand2_1
XANTENNA__12107__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13275_ clknet_leaf_153_clk _00506_ net1117 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[263\]
+ sky130_fd_sc_hd__dfrtp_1
X_12226_ net592 _06154_ net518 net379 net1653 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__a32o_1
XANTENNA__12191__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08934__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ net184 net2405 net387 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__mux2_1
XANTENNA__06945__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11108_ _05818_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__xnor2_1
X_12088_ net589 _06053_ net516 net394 net1693 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__a32o_1
XANTENNA__08320__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11039_ _05761_ _05762_ _05737_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_34_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07444__B _02394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12494__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06580_ final_design.cpu.reg_window\[605\] final_design.cpu.reg_window\[637\] net957
+ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__mux2_1
XANTENNA__09647__B1 _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08250_ final_design.cpu.reg_window\[330\] final_design.cpu.reg_window\[362\] net839
+ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__mux2_1
XANTENNA__09662__A3 _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08870__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07201_ final_design.cpu.reg_window\[649\] final_design.cpu.reg_window\[681\] net924
+ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08181_ net604 _03129_ _03105_ _01966_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__o211a_1
XFILLER_0_172_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07132_ final_design.cpu.reg_window\[907\] final_design.cpu.reg_window\[939\] net945
+ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07063_ net768 _02013_ net754 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08230__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ _02912_ _02913_ _02914_ _02915_ net683 net705 vssd1 vssd1 vccd1 vccd1 _02916_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout382_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _04116_ _04310_ _04621_ net498 _04622_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__a221oi_4
X_06916_ _01863_ _01864_ _01865_ _01866_ net774 net795 vssd1 vssd1 vccd1 vccd1 _01867_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07036__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12485__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07896_ final_design.cpu.reg_window\[215\] final_design.cpu.reg_window\[247\] net843
+ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__mux2_1
XANTENNA__09850__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09635_ _03031_ _04430_ _02997_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__o21ai_1
X_06847_ final_design.cpu.reg_window\[20\] final_design.cpu.reg_window\[52\] net947
+ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07361__A1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout268_X net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06778_ final_design.cpu.reg_window\[406\] final_design.cpu.reg_window\[438\] net902
+ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__mux2_1
XANTENNA__06685__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ net549 net548 net547 net546 net453 net462 vssd1 vssd1 vccd1 vccd1 _04485_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08466__A _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11445__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08517_ net729 _03467_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07113__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09497_ net473 _04086_ _04411_ _04415_ _04410_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__o311a_1
XFILLER_0_136_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07113__B2 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1177_X net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08448_ final_design.cpu.reg_window\[196\] final_design.cpu.reg_window\[228\] net858
+ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08379_ final_design.cpu.reg_window\[390\] final_design.cpu.reg_window\[422\] net831
+ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10410_ _03352_ _05181_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11390_ net437 net593 _06075_ net318 net1750 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__a32o_1
XANTENNA__06624__A0 final_design.cpu.reg_window\[411\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10341_ net1595 net1024 net1001 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1
+ vccd1 _00098_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10420__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13060_ clknet_leaf_107_clk _00291_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_10272_ _05133_ net809 _05132_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout971_X net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12011_ _06213_ net280 net400 net2327 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__a22o_1
XANTENNA__11766__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11993__C net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 net461 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__clkbuf_4
Xfanout471 net473 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_4
Xfanout482 _03484_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13962_ clknet_leaf_3_clk _01193_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[950\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout493 net495 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12476__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ clknet_leaf_90_clk _00151_ net1232 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11684__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ clknet_leaf_149_clk _01124_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[881\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07551__Y _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12844_ clknet_leaf_86_clk _00082_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11726_ net593 net424 _06221_ net298 net1867 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__a32o_1
XFILLER_0_166_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06863__B1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11657_ net187 net640 vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10608_ _05349_ _05350_ _05331_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12400__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08315__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11588_ net188 net644 vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold908 final_design.cpu.reg_window\[513\] vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13327_ clknet_leaf_90_clk _00558_ net1232 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[315\]
+ sky130_fd_sc_hd__dfrtp_1
X_10539_ net1583 net1045 net1017 _05286_ vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__a22o_1
Xhold919 final_design.cpu.reg_window\[929\] vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13258_ clknet_leaf_0_clk _00489_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[246\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12209_ net579 _06137_ net511 net377 net1664 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__a32o_1
X_13189_ clknet_leaf_5_clk _00420_ net1096 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[177\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07455__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08050__S net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07750_ net621 _02698_ _02699_ net559 vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12467__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06701_ final_design.cpu.reg_window\[665\] final_design.cpu.reg_window\[697\] net940
+ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07681_ final_design.cpu.reg_window\[542\] final_design.cpu.reg_window\[574\] net850
+ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__mux2_1
XANTENNA__07343__B2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09420_ net485 _04338_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__nand2_1
X_06632_ net765 _01576_ net757 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__o21a_1
XANTENNA__12300__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07190__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06563_ final_design.cpu.reg_window\[413\] final_design.cpu.reg_window\[445\] net962
+ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__mux2_1
X_09351_ _02671_ _04094_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08302_ final_design.cpu.reg_window\[969\] final_design.cpu.reg_window\[1001\] net842
+ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09282_ net549 net548 net547 net546 net457 net467 vssd1 vssd1 vccd1 vccd1 _04201_
+ sky130_fd_sc_hd__mux4_1
X_06494_ net760 _01444_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ final_design.cpu.reg_window\[907\] final_design.cpu.reg_window\[939\] net857
+ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout228_A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ _03111_ _03112_ _03113_ _03114_ net683 net705 vssd1 vssd1 vccd1 vccd1 _03115_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09399__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08225__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07115_ _02058_ _02063_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08095_ _03042_ _03043_ _03044_ _03045_ net687 net708 vssd1 vssd1 vccd1 vccd1 _03046_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload70 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__inv_6
XANTENNA_fanout1137_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07046_ net1053 _01409_ net1003 final_design.reqhand.instruction\[14\] vssd1 vssd1
+ vccd1 vccd1 _01997_ sky130_fd_sc_hd__a31o_1
Xclkload81 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload92 clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 clkload92/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_149_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout597_A _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07031__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08997_ _03738_ _03739_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__A0 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ net608 _02894_ _02869_ _01750_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_3_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11666__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ net891 _02811_ _02817_ _02823_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__o32a_4
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09618_ _04059_ net321 vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10890_ net49 _05620_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__xor2_1
XANTENNA__08196__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09549_ _04342_ _04460_ _04465_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_167_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12091__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12560_ _06223_ net359 net326 net2414 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11511_ net2242 net217 net525 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12491_ _06151_ net356 net333 net2399 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14230_ net1295 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_110_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11442_ net817 _02359_ _02392_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12394__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11197__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14161_ clknet_leaf_82_clk _01335_ net1247 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11373_ net658 net184 vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_169_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input60_A mem_adr_start[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10324_ net1505 net1024 net1001 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1
+ vccd1 _00081_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13112_ clknet_leaf_133_clk _00343_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14092_ clknet_leaf_71_clk _01289_ net1243 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11496__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10255_ final_design.uart.BAUD_counter\[19\] final_design.uart.BAUD_counter\[20\]
+ _05119_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13043_ clknet_leaf_33_clk _00274_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08445__S0 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1200 net1217 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__clkbuf_4
Xfanout1211 net1216 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12889__Q final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ final_design.uart.BAUD_counter\[13\] final_design.uart.BAUD_counter\[12\]
+ final_design.uart.BAUD_counter\[15\] final_design.uart.BAUD_counter\[14\] vssd1
+ vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__or4_1
Xfanout1222 net1223 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1233 net1234 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__buf_2
Xfanout1244 net1246 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__clkbuf_4
Xfanout1255 net1256 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__buf_2
Xfanout290 net294 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07562__X _02513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09314__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13945_ clknet_leaf_165_clk _01176_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[933\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12120__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13876_ clknet_leaf_103_clk _01107_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[864\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09078__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12827_ net1357 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12779__10 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__inv_2
XANTENNA__12082__B1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12758_ _06383_ _06390_ _06391_ _06333_ final_design.VGA_adr\[6\] vssd1 vssd1 vccd1
+ vccd1 _06395_ sky130_fd_sc_hd__a32o_1
XANTENNA__08834__A final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07184__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11709_ net199 net634 vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__and2_1
XANTENNA__10575__S net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12689_ _01401_ _05038_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold705 final_design.cpu.reg_window\[856\] vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold716 final_design.cpu.reg_window\[1018\] vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 final_design.cpu.reg_window\[434\] vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 final_design.cpu.reg_window\[534\] vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold749 final_design.cpu.reg_window\[386\] vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11259__X _05960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08920_ final_design.CPU_instr_adr\[22\] _01756_ _03862_ vssd1 vssd1 vccd1 vccd1
+ _03863_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11345__C1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11896__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09952__X _04871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ final_design.CPU_instr_adr\[30\] _03801_ vssd1 vssd1 vccd1 vccd1 _03802_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07802_ final_design.cpu.reg_window\[793\] final_design.cpu.reg_window\[825\] net866
+ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__mux2_1
X_08782_ _03688_ _03732_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_58_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08568__X _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07472__X _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11648__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ _02680_ _02681_ _02682_ _02683_ net695 net713 vssd1 vssd1 vccd1 vccd1 _02684_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_140_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout178_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12030__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ final_design.cpu.reg_window\[414\] final_design.cpu.reg_window\[446\] net849
+ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09403_ _02576_ _02606_ _04171_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06615_ net898 _01559_ _01565_ _01547_ _01553_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__a32oi_4
X_07595_ _01539_ net613 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__nand2_1
XANTENNA__13423__Q final_design.cpu.reg_window\[411\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09334_ _04249_ _04251_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__xnor2_1
X_06546_ _01485_ _01489_ net741 _01495_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__and4_2
XFILLER_0_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12073__B1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08277__C1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10623__A1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11820__A0 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09265_ net71 _04183_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__or2_1
X_12778__9 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__inv_2
X_06477_ final_design.cpu.reg_window\[478\] final_design.cpu.reg_window\[510\] net930
+ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout512_A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1254_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11170__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06922__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08216_ _03103_ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__nand2_1
X_09196_ _02545_ _04088_ _04096_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12376__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11179__A2 _05143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13755__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout300_X net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08147_ _02030_ net616 vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08044__A2 _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07794__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09575__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09792__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ _03028_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout881_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07029_ _01976_ _01977_ _01978_ _01979_ net780 net792 vssd1 vssd1 vccd1 vccd1 _01980_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_112_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap980 _01472_ vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ _04637_ _04924_ _04958_ _04574_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__and4b_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11887__A0 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold10 final_design.cpu.reg_window\[30\] vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 final_design.cpu.reg_window\[12\] vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 net104 vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 final_design.cpu.reg_window\[6\] vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 final_design.cpu.reg_window\[5\] vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 final_design.VGA_data_control.data_to_VGA\[27\] vssd1 vssd1 vccd1 vccd1 net1418
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 final_design.VGA_data_control.data_to_VGA\[13\] vssd1 vssd1 vccd1 vccd1 net1429
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 net165 vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 final_design.cpu.reg_window\[11\] vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ net230 net2382 net402 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__mux2_1
XANTENNA__12300__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13730_ clknet_leaf_28_clk _00961_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[718\]
+ sky130_fd_sc_hd__dfrtp_1
X_10942_ _05646_ _05667_ net243 vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_168_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07034__S net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13661_ clknet_leaf_11_clk _00892_ net1129 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[649\]
+ sky130_fd_sc_hd__dfrtp_1
X_10873_ _05508_ _05542_ _05603_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__o31a_1
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12612_ net1425 net1009 net995 final_design.data_from_mem\[30\] vssd1 vssd1 vccd1
+ vccd1 _01305_ sky130_fd_sc_hd__a22o_1
XANTENNA__07969__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12064__B1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13592_ clknet_leaf_131_clk _00823_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[580\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08654__A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12543_ _06206_ net349 net324 net1588 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09480__A1 _04398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12474_ _06134_ net351 net332 net2420 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12367__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10408__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ net1282 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_124_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11425_ net2002 net205 net311 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14144_ clknet_leaf_77_clk _01318_ net1253 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11356_ net657 net189 vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10307_ _01384_ net1061 _05160_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__or3b_1
X_14075_ clknet_leaf_52_clk _01272_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12115__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11287_ net669 _03912_ net743 vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a21o_1
XANTENNA__07209__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13026_ clknet_leaf_27_clk _00257_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10238_ final_design.uart.BAUD_counter\[13\] final_design.uart.BAUD_counter\[12\]
+ _05108_ final_design.uart.BAUD_counter\[14\] vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__a31o_1
XANTENNA__11878__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1030 _01411_ vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_4
Xfanout1041 net1043 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__buf_2
X_10169_ final_design.vga.h_current_state\[0\] final_design.vga.h_current_state\[1\]
+ _05044_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__o21ai_1
Xfanout1052 _01394_ vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__buf_1
Xfanout1063 final_design.VGA_data_control.h_count\[1\] vssd1 vssd1 vccd1 vccd1 net1063
+ sky130_fd_sc_hd__buf_4
Xfanout1074 net1075 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1085 net1104 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_4
Xfanout1096 net1099 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_4
X_13928_ clknet_leaf_120_clk _01159_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[916\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_164_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07849__A2 _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10853__A1 _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13859_ clknet_leaf_5_clk _01090_ net1096 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[847\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06521__A2 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11542__X _06127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07380_ _02326_ _02330_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__nand2_1
XANTENNA__06783__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08564__A _02394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11802__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09471__A1 _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09050_ _02442_ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08001_ final_design.cpu.reg_window\[976\] final_design.cpu.reg_window\[1008\] net878
+ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold502 final_design.cpu.reg_window\[603\] vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold513 final_design.cpu.reg_window\[590\] vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold524 final_design.cpu.reg_window\[744\] vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold535 final_design.cpu.reg_window\[896\] vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06588__A2 _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold546 final_design.cpu.reg_window\[209\] vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold557 final_design.cpu.reg_window\[348\] vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 final_design.cpu.reg_window\[779\] vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11581__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold579 final_design.cpu.reg_window\[344\] vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ net496 _04868_ _04869_ _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08903_ _01661_ _01662_ _02469_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__or3_1
XANTENNA__07119__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11869__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ _04341_ _04801_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__or2_1
XANTENNA__11333__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 final_design.CPU_instr_adr\[7\] vssd1 vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ final_design.CPU_instr_adr\[5\] _03784_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__and2_1
Xhold1213 final_design.VGA_adr\[9\] vssd1 vssd1 vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1002_A _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10988__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ final_design.CPU_instr_adr\[1\] _02391_ _02393_ vssd1 vssd1 vccd1 vccd1 _03716_
+ sky130_fd_sc_hd__nand3b_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07716_ net723 _02666_ net893 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12294__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08696_ _01487_ _03646_ _02094_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_68_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout250_X net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07647_ final_design.cpu.reg_window\[604\] final_design.cpu.reg_window\[636\] net871
+ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout727_A _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07789__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07578_ final_design.cpu.reg_window\[543\] final_design.cpu.reg_window\[575\] net846
+ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12597__B2 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__Y _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09317_ net480 _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__nor2_1
X_06529_ _01478_ _01479_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_118_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ _04158_ _04164_ _04166_ _04133_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09179_ net530 net468 net459 vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__or3_1
XANTENNA__11021__A1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ _03620_ _05854_ _05906_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__and3_2
XFILLER_0_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12190_ net1679 net186 net382 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout884_X net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11141_ final_design.reqhand.data_from_UART\[0\] final_design.data_from_mem\[0\]
+ net249 vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07871__S1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11072_ _05773_ _05791_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__and2_1
Xinput100 nrst vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__buf_4
X_10023_ net68 _04940_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__or2_1
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12285__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ _06176_ net293 net407 net1570 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__a22o_1
X_13713_ clknet_leaf_107_clk _00944_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[701\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10925_ _05652_ _05653_ _05632_ _05634_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_169_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13644_ clknet_leaf_125_clk _00875_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[632\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10856_ net80 net1055 vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12588__B2 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13575_ clknet_leaf_8_clk _00806_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[563\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09453__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ net43 _05521_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11260__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12526_ _06188_ net357 net329 net2111 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10853__S net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12457_ net2141 net189 net337 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11408_ net817 _02359_ net815 vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_10_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12388_ net2058 net191 net272 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11563__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06931__A_N net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14127_ clknet_leaf_75_clk final_design.vga.v_next_count\[7\] net1245 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[7\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_91_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11339_ _06027_ _06029_ _06030_ net598 vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__o211a_2
XFILLER_0_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14058_ clknet_leaf_46_clk _00020_ net1148 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11315__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ net1351 _00240_ net1224 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__06778__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06880_ net759 _01830_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__nor2_1
XANTENNA__11256__Y _05958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12276__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08550_ final_design.cpu.reg_window\[833\] final_design.cpu.reg_window\[865\] net854
+ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__mux2_1
XANTENNA__09141__A0 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07501_ _02002_ _02450_ _02001_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08481_ final_design.cpu.reg_window\[67\] final_design.cpu.reg_window\[99\] net864
+ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12291__A3 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11713__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07432_ final_design.cpu.reg_window\[705\] final_design.cpu.reg_window\[737\] net932
+ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06807__A _01750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07402__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07363_ final_design.cpu.reg_window\[771\] final_design.cpu.reg_window\[803\] net944
+ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06526__B _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09102_ _02364_ _02429_ net628 vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10054__A2 _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11251__A1 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07294_ final_design.cpu.reg_window\[197\] final_design.cpu.reg_window\[229\] net904
+ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09033_ final_design.CPU_instr_adr\[11\] _03788_ vssd1 vssd1 vccd1 vccd1 _03964_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_A _05958_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout308_A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07638__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12200__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 final_design.cpu.reg_window\[521\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__C1 _02239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08233__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold321 final_design.cpu.reg_window\[956\] vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 final_design.cpu.reg_window\[862\] vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07302__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 final_design.cpu.reg_window\[655\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 final_design.cpu.reg_window\[185\] vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold365 final_design.cpu.reg_window\[216\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 final_design.VGA_data_control.ready_data\[7\] vssd1 vssd1 vccd1 vccd1 net1729
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1217_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 final_design.cpu.reg_window\[131\] vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout801 net807 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__buf_2
Xhold398 final_design.cpu.reg_window\[600\] vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout812 _05090_ vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_2
X_09935_ net491 _04619_ _04852_ _04853_ _04341_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a221o_1
XANTENNA__12982__RESET_B net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout823 net829 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_2
Xfanout834 net835 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout677_A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__A2 _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net855 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_2
Xfanout856 net857 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__clkbuf_4
Xfanout867 net876 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_2
XANTENNA__06688__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09866_ _03294_ _03568_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__xnor2_1
Xhold1010 final_design.cpu.reg_window\[741\] vssd1 vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07605__S1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout878 net886 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_4
Xhold1021 final_design.cpu.reg_window\[495\] vssd1 vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09380__A0 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07373__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout889 net890 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_8
X_08817_ _03753_ _03763_ _03767_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__o21ba_1
Xhold1032 final_design.cpu.reg_window\[547\] vssd1 vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 final_design.cpu.reg_window\[555\] vssd1 vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1054 final_design.cpu.reg_window\[343\] vssd1 vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _03358_ net447 _04242_ _04086_ _04715_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout844_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 final_design.cpu.reg_window\[932\] vssd1 vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1076 final_design.cpu.reg_window\[324\] vssd1 vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ _03697_ _03698_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12267__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1087 final_design.cpu.reg_window\[810\] vssd1 vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 final_design.cpu.reg_window\[633\] vssd1 vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_159_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ _03629_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__inv_2
XANTENNA__12282__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10710_ _05447_ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__nand2_1
XANTENNA__12019__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11690_ net429 net577 _06203_ net296 net1852 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__a32o_1
XANTENNA__06717__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13770__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10641_ _05347_ _05364_ _05383_ _05362_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13360_ clknet_leaf_112_clk _00591_ net1212 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[348\]
+ sky130_fd_sc_hd__dfrtp_1
X_10572_ _05291_ _05294_ _05316_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11793__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11769__S net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12311_ net1590 net207 net365 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13291_ clknet_leaf_21_clk _00522_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[279\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09738__A2 _04639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12242_ net579 _06172_ net511 net373 net1434 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__a32o_1
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11545__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ net1792 net217 net381 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__mux2_1
XANTENNA__07844__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124_ net679 _02358_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__or3_4
X_11055_ _04325_ net249 net678 vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06598__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ _04614_ _04615_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__nor2_1
XANTENNA__12897__Q final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09910__A2 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12258__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08666__X _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ net433 net565 net640 vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__and3_1
XFILLER_0_157_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12273__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06488__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ net972 _05636_ _05637_ net968 vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08318__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11888_ net227 net1952 net276 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13627_ clknet_leaf_156_clk _00858_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[615\]
+ sky130_fd_sc_hd__dfrtp_1
X_10839_ _05570_ _05571_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__xor2_1
XFILLER_0_116_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8__f_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_41_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11233__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ clknet_leaf_130_clk _00789_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[546\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ _06171_ net353 net329 net1822 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13489_ clknet_leaf_108_clk _00720_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[477\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09729__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10744__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07892__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07981_ net609 _02929_ _02905_ net548 vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__o211a_2
XFILLER_0_38_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11267__X _05967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ _04627_ _04638_ net448 vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__a21o_1
X_06932_ net550 _01881_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__xor2_1
XANTENNA__12303__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ net448 _04569_ _04566_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__o21a_1
X_06863_ net772 _01813_ net898 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08260__S1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ net614 _03550_ _03524_ _02419_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__o211a_1
XANTENNA__07912__B2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12249__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09582_ _03582_ _04499_ _03134_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__a21oi_1
X_06794_ final_design.cpu.reg_window\[790\] final_design.cpu.reg_window\[822\] net905
+ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08533_ net622 _03481_ _03482_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_65_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08468__A2 _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08736__B _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08464_ _03402_ _03403_ _03414_ net892 vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_102_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07132__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07415_ final_design.cpu.reg_window\[257\] final_design.cpu.reg_window\[289\] net930
+ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09417__A1 _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ final_design.cpu.reg_window\[710\] final_design.cpu.reg_window\[742\] net830
+ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout425_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1167_A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11224__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07346_ net752 net675 net731 _01496_ _02296_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__o221a_2
XANTENNA__12421__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09848__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08752__A final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11775__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07277_ final_design.cpu.reg_window\[838\] final_design.cpu.reg_window\[870\] net913
+ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09016_ final_design.CPU_instr_adr\[12\] _03789_ final_design.CPU_instr_adr\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout794_A _01419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08928__B1 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold140 final_design.VGA_data_control.ready_data\[30\] vssd1 vssd1 vccd1 vccd1 net1493
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold151 final_design.cpu.reg_window\[972\] vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 final_design.cpu.reg_window\[522\] vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 final_design.cpu.reg_window\[458\] vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 final_design.cpu.reg_window\[528\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 final_design.VGA_data_control.ready_data\[18\] vssd1 vssd1 vccd1 vccd1 net1548
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout961_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout620 _02513_ vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_2
Xfanout631 _02506_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_2
Xfanout642 _06123_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_4
XANTENNA__07374__Y _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09918_ net486 _04407_ _04835_ _04219_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_109_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout653 _05853_ vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12488__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout664 _05142_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_4
Xfanout675 _01498_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_2
Xfanout686 net698 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_8
X_09849_ _04751_ _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout697 net698 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__buf_4
XANTENNA__11160__B1 _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ clknet_leaf_79_clk _00098_ net1250 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11811_ net231 net2284 net268 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__mux2_1
XANTENNA__08003__S1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12255__A3 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11742_ net238 net2337 net417 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11673_ net228 net635 vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07977__S net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13412_ clknet_leaf_100_clk _00643_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[400\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10018__A2 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input90_A memory_size[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ _04745_ net247 net678 vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_12_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12412__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06881__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13343_ clknet_leaf_136_clk _00574_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[331\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10555_ net63 _05301_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13274_ clknet_leaf_151_clk _00505_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[262\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ net90 final_design.VGA_adr\[0\] vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12225_ net590 _06153_ net516 net378 net1612 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__a32o_1
XFILLER_0_102_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12156_ net186 net2352 net387 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11107_ net60 _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12123__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12479__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12087_ net585 _06046_ net517 net394 net2078 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_142_Left_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11038_ net88 net1058 vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09647__A1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12989_ net1331 _00220_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_151_Left_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07200_ final_design.cpu.reg_window\[713\] final_design.cpu.reg_window\[745\] net924
+ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12403__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08180_ _01967_ net616 vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07131_ final_design.cpu.reg_window\[971\] final_design.cpu.reg_window\[1003\] net938
+ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__mux2_1
XANTENNA__08622__A2 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07062_ _02009_ _02010_ _02011_ _02012_ net777 net797 vssd1 vssd1 vccd1 vccd1 _02013_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_4__f_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_160_Left_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12033__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ final_design.cpu.reg_window\[145\] final_design.cpu.reg_window\[177\] net827
+ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09703_ net490 _04578_ _04579_ _04620_ _04341_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_96_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06915_ final_design.cpu.reg_window\[146\] final_design.cpu.reg_window\[178\] net901
+ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07895_ final_design.cpu.reg_window\[23\] final_design.cpu.reg_window\[55\] net843
+ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__mux2_1
XANTENNA__09886__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09886__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09634_ _02997_ _03031_ _04430_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__or3_1
X_06846_ final_design.cpu.reg_window\[84\] final_design.cpu.reg_window\[116\] net949
+ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09565_ _03134_ _04087_ _04483_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__a21oi_1
X_06777_ final_design.cpu.reg_window\[470\] final_design.cpu.reg_window\[502\] net903
+ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout542_A _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12237__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08516_ _03463_ _03464_ _03465_ _03466_ net693 net712 vssd1 vssd1 vccd1 vccd1 _03467_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_121_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09496_ net481 _04086_ _04412_ _04414_ _04269_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__o311a_1
XANTENNA__07113__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08310__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11996__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08447_ final_design.cpu.reg_window\[4\] final_design.cpu.reg_window\[36\] net858
+ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_171_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_171_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1072_X net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_A _01418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07797__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06554__X _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08378_ final_design.cpu.reg_window\[454\] final_design.cpu.reg_window\[486\] net835
+ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07329_ _02276_ _02277_ _02278_ _02279_ net783 net802 vssd1 vssd1 vccd1 vccd1 _02280_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_104_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10340_ net1531 net1025 net1002 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1
+ vccd1 _00097_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10420__A2 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10271_ final_design.uart.BAUD_counter\[25\] final_design.uart.BAUD_counter\[26\]
+ _05129_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__and3_1
X_12010_ _06212_ net278 net400 net2161 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11348__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout450 _04070_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_4
Xfanout461 _03551_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_2
Xfanout472 net473 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__dlymetal6s2s_1
X_13961_ clknet_leaf_88_clk _01192_ net1235 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[949\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09877__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout483 net489 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__buf_2
Xfanout494 net495 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_2
X_12912_ clknet_leaf_33_clk _00150_ net1130 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09760__B _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11684__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13892_ clknet_leaf_100_clk _01123_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[880\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07561__A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ clknet_leaf_86_clk _00081_ net1249 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12228__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11083__A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11436__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_15__f_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11987__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11725_ net185 net637 vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_162_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_162_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input93_X net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06863__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11656_ net435 net591 _06185_ net301 net1610 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__a32o_1
XFILLER_0_154_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06905__A _01850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10607_ _05331_ _05349_ _05350_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__and3b_1
X_11587_ net434 net586 _06149_ net305 net1617 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12118__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13326_ clknet_leaf_113_clk _00557_ net1212 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[314\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06615__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10538_ _05268_ _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__xnor2_1
Xhold909 final_design.cpu.reg_window\[950\] vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13257_ clknet_leaf_85_clk _00488_ net1235 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[245\]
+ sky130_fd_sc_hd__dfrtp_1
X_10469_ net36 _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12208_ net584 _06136_ net514 net378 net1994 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_36_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08331__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13188_ clknet_leaf_94_clk _00419_ net1227 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[176\]
+ sky130_fd_sc_hd__dfrtp_1
X_12139_ net217 net2514 net385 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07591__A2 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06700_ final_design.cpu.reg_window\[729\] final_design.cpu.reg_window\[761\] net940
+ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07680_ final_design.cpu.reg_window\[606\] final_design.cpu.reg_window\[638\] net850
+ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06631_ net773 _01581_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__or2_1
XANTENNA__11705__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12219__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09350_ net496 _04268_ _04231_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a21o_1
X_06562_ final_design.cpu.reg_window\[477\] final_design.cpu.reg_window\[509\] net962
+ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08301_ final_design.cpu.reg_window\[777\] final_design.cpu.reg_window\[809\] net843
+ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__mux2_1
XANTENNA__11978__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09281_ net554 net553 net552 net551 net458 net466 vssd1 vssd1 vccd1 vccd1 _04200_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06493_ _01440_ _01441_ _01442_ _01443_ net781 net799 vssd1 vssd1 vccd1 vccd1 _01444_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_153_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_153_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08573__Y _03524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11280__X _05979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08232_ final_design.cpu.reg_window\[971\] final_design.cpu.reg_window\[1003\] net877
+ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__mux2_1
XANTENNA__11721__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08163_ final_design.cpu.reg_window\[143\] final_design.cpu.reg_window\[175\] net824
+ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12028__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__B1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07114_ _02059_ _02064_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_166_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ final_design.cpu.reg_window\[396\] final_design.cpu.reg_window\[428\] net846
+ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload60 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__clkinv_2
Xclkload71 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_77_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07045_ net896 _01988_ _01994_ _01981_ _01982_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a32o_2
XFILLER_0_113_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload82 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 clkload82/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_149_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload93 clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_149_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09020__A2 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout492_A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07031__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10072__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ net257 _03930_ net1026 vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_145_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ net554 _02896_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout280_X net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11666__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06696__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ net729 _02828_ net891 vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_173_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07381__A _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07965__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _04066_ _04108_ net319 vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__o21ai_1
X_06829_ final_design.cpu.reg_window\[597\] final_design.cpu.reg_window\[629\] net963
+ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__mux2_1
XANTENNA__11615__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout924_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11418__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09548_ net320 _04373_ _04376_ net321 _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11969__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12091__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_144_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_144_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09479_ _04396_ _04397_ net480 vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__mux2_2
XFILLER_0_148_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11631__A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ net2126 net219 net524 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12490_ _06150_ net353 net333 net2208 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07320__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11441_ net1614 net176 net312 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08598__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14160_ clknet_leaf_80_clk _01334_ net1248 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11372_ net599 _06058_ _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__and3_2
XFILLER_0_116_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13111_ clknet_leaf_145_clk _00342_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10323_ net1586 net1024 net1001 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1
+ vccd1 _00080_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14091_ clknet_leaf_71_clk _01288_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input53_A mem_adr_start[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ clknet_leaf_44_clk _00273_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10254_ final_design.uart.BAUD_counter\[19\] final_design.uart.BAUD_counter\[18\]
+ _05118_ final_design.uart.BAUD_counter\[20\] vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__a31o_1
XANTENNA__11354__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08445__S1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__clkbuf_4
Xfanout1212 net1216 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__clkbuf_4
Xfanout1223 net1224 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_2
X_10185_ final_design.uart.BAUD_counter\[9\] final_design.uart.BAUD_counter\[8\] final_design.uart.BAUD_counter\[11\]
+ final_design.uart.BAUD_counter\[10\] vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__or4b_1
XANTENNA__11087__A1_N net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07990__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1234 net1239 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__buf_2
Xfanout1245 net1246 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_4
Xfanout1256 net100 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout280 net283 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_4
Xfanout291 net294 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13284__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__A3 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13944_ clknet_leaf_138_clk _01175_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[932\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07291__A _02239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13875_ clknet_leaf_30_clk _01106_ net1139 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[863\]
+ sky130_fd_sc_hd__dfrtp_1
X_12826_ net1366 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10880__A2 _05610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12757_ _06392_ _06393_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__or2_1
XANTENNA__12196__X _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08825__A2 _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_135_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_167_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07184__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06836__A1 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ net566 net420 _06212_ net295 net1973 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12688_ _06331_ net1420 net991 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08326__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11639_ net203 net638 vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__and2_1
X_12794__25 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__inv_2
XFILLER_0_13_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold706 final_design.cpu.reg_window\[739\] vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11593__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 final_design.cpu.reg_window\[321\] vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold728 final_design.cpu.reg_window\[413\] vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ clknet_leaf_30_clk _00540_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[297\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold739 final_design.uart.working_data\[7\] vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09538__A0 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09002__A2 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11345__B1 _06035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10604__B _04787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08850_ final_design.CPU_instr_adr\[29\] _03800_ vssd1 vssd1 vccd1 vccd1 _03801_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07801_ final_design.cpu.reg_window\[857\] final_design.cpu.reg_window\[889\] net866
+ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__mux2_1
X_08781_ _03692_ _03694_ _03729_ _03690_ _03689_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__a311o_1
XFILLER_0_58_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11648__A1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ final_design.cpu.reg_window\[154\] final_design.cpu.reg_window\[186\] net872
+ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__mux2_1
XANTENNA__12311__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__B _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09710__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ final_design.cpu.reg_window\[478\] final_design.cpu.reg_window\[510\] net849
+ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__mux2_1
XANTENNA__10320__B2 final_design.data_from_mem\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09402_ _04051_ _04291_ _04292_ _04320_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__o31a_1
XFILLER_0_153_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06614_ net771 _01564_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__or2_1
XANTENNA__09069__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07594_ _02543_ _02544_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__or2_2
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09333_ _04251_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06545_ _01489_ net741 _01495_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__and3_1
XANTENNA__12936__RESET_B net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_A _05890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_126_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_164_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08744__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout338_A _06282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ net69 _04182_ net70 vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06476_ final_design.data_from_mem\[18\] net981 _01425_ vssd1 vssd1 vccd1 vccd1 _01427_
+ sky130_fd_sc_hd__o21ai_2
XANTENNA__08236__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06922__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08215_ _03132_ _03133_ _03162_ _03163_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09195_ _02543_ net445 _04113_ net530 vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout505_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08146_ net605 _03096_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06686__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08077_ _03025_ _03027_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__nor2_2
XANTENNA__09792__A3 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09529__B1 _04231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07376__A final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07028_ final_design.cpu.reg_window\[14\] final_design.cpu.reg_window\[46\] net926
+ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold11 final_design.cpu.reg_window\[8\] vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09591__A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 final_design.cpu.reg_window\[22\] vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 final_design.cpu.reg_window\[2\] vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 final_design.VGA_data_control.data_to_VGA\[11\] vssd1 vssd1 vccd1 vccd1 net1397
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ net630 _03914_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__a21o_1
Xhold55 final_design.cpu.reg_window\[15\] vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 net137 vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 net145 vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 net139 vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11990_ net681 _06118_ _06193_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__or3_1
Xhold99 final_design.cpu.reg_window\[960\] vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_168_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10941_ _05662_ _05643_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout927_X net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13660_ clknet_leaf_152_clk _00891_ net1117 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[648\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10872_ _05560_ _05578_ _05603_ _05563_ _05580_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12611_ net1632 net1011 net997 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1
+ vccd1 _01304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13591_ clknet_leaf_136_clk _00822_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[579\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_117_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08363__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12542_ _06205_ net353 net325 net2170 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11080__B net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ _06133_ net348 net332 net2088 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14212_ net1281 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_149_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11424_ net1676 net207 net312 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__mux2_1
XANTENNA__10378__B2 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ clknet_leaf_75_clk _01317_ net1253 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11355_ _06041_ _06043_ _06044_ net599 vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__o211a_2
XFILLER_0_1_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10306_ final_design.VGA_data_control.data_to_VGA\[27\] final_design.VGA_data_control.data_to_VGA\[26\]
+ final_design.VGA_data_control.data_to_VGA\[25\] final_design.VGA_data_control.data_to_VGA\[24\]
+ net1063 net1062 vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__mux4_1
X_14074_ clknet_leaf_53_clk _01271_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11286_ final_design.data_from_mem\[17\] net235 net233 vssd1 vssd1 vccd1 vccd1 _05984_
+ sky130_fd_sc_hd__a21o_2
XANTENNA__14180__Q final_design.VGA_adr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13025_ clknet_leaf_159_clk _00256_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10237_ net1539 _05109_ _05111_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__a21oi_1
Xfanout1020 _05171_ vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_4
Xfanout1031 final_design.CPU_instr_adr\[2\] vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_4
Xfanout1042 net1044 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__dlymetal6s2s_1
X_14193__1321 vssd1 vssd1 vccd1 vccd1 net1321 _14193__1321/LO sky130_fd_sc_hd__conb_1
XANTENNA__09940__B1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10168_ _05041_ _05060_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[8\]
+ sky130_fd_sc_hd__nor2_1
Xfanout1053 _01393_ vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__buf_2
Xfanout1064 final_design.VGA_data_control.v_count\[4\] vssd1 vssd1 vccd1 vccd1 net1064
+ sky130_fd_sc_hd__buf_2
XANTENNA__08829__B _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1075 net1080 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_4
Xfanout1086 net1104 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12131__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1097 net1099 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10440__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10099_ _05011_ _05014_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__or2_1
XANTENNA__07929__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13927_ clknet_leaf_13_clk _01158_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[915\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06601__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13858_ clknet_leaf_14_clk _01089_ net1103 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[846\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12809_ net1392 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12055__A1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_108_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13789_ clknet_leaf_13_clk _01020_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[777\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08000_ final_design.cpu.reg_window\[784\] final_design.cpu.reg_window\[816\] net878
+ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12358__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10369__B2 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07234__A1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold503 final_design.cpu.reg_window\[797\] vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold514 final_design.cpu.reg_window\[251\] vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 final_design.cpu.reg_window\[332\] vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12306__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10615__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold536 final_design.cpu.reg_window\[687\] vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold547 final_design.cpu.reg_window\[1000\] vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07785__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold558 final_design.cpu.reg_window\[477\] vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _04091_ _04436_ _04446_ net496 vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a31oi_1
Xhold569 final_design.cpu.reg_window\[503\] vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
X_08902_ _03771_ _03846_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_70_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09882_ net487 _04733_ _04799_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__o22a_1
X_08833_ final_design.CPU_instr_adr\[4\] final_design.CPU_instr_adr\[3\] net1031 vssd1
+ vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__and3_1
XANTENNA__07924__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1203 net117 vssd1 vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 final_design.VGA_adr\[2\] vssd1 vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout190_A _06038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__B _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout288_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ final_design.CPU_instr_adr\[0\] _02425_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__and2_1
XANTENNA__12041__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07135__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07715_ _02662_ _02663_ _02664_ _02665_ net697 net715 vssd1 vssd1 vccd1 vccd1 _02666_
+ sky130_fd_sc_hd__mux4_1
X_08695_ _01998_ _02028_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout455_A net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1197_A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07646_ final_design.cpu.reg_window\[668\] final_design.cpu.reg_window\[700\] net871
+ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10349__X _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07577_ final_design.cpu.reg_window\[607\] final_design.cpu.reg_window\[639\] net846
+ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__mux2_1
XANTENNA__10057__B1 _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ net536 net534 net533 _02325_ net460 net470 vssd1 vssd1 vccd1 vccd1 _04235_
+ sky130_fd_sc_hd__mux4_1
X_06528_ _01393_ net1006 net1003 _01378_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__a31o_1
XANTENNA__11254__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07473__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09247_ _02673_ _02705_ _02738_ _02770_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06459_ net1068 net1050 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12349__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13976__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09178_ net494 _03629_ net666 vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__or3_4
XFILLER_0_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11557__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08129_ final_design.cpu.reg_window\[205\] final_design.cpu.reg_window\[237\] net830
+ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__mux2_1
X_11140_ net653 _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__and2_2
XFILLER_0_102_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11309__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ _05757_ _05775_ _05792_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__or3_1
X_10022_ net68 _04940_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__nand2_1
XANTENNA__12521__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__B2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06831__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12285__A1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _06175_ net280 net404 net1737 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__a22o_1
X_10924_ net82 net1060 net83 vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__or3b_1
X_13712_ clknet_leaf_105_clk _00943_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[700\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06884__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08665__A _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10855_ _05549_ _05570_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__nor2_1
X_13643_ clknet_leaf_16_clk _00874_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[631\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11245__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13574_ clknet_leaf_169_clk _00805_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[562\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ net43 _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09453__A2 _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10419__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12525_ _06187_ net358 net329 net2027 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12456_ net2411 net191 net337 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ net428 net580 _06090_ net316 net1552 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_10_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12126__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12387_ net1651 net193 net270 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14126_ clknet_leaf_75_clk final_design.vga.v_next_count\[6\] net1252 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[6\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_91_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11338_ _04546_ _04549_ net659 vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_91_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14057_ clknet_leaf_47_clk _00019_ net1148 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11269_ net744 _03930_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13008_ net1350 _00239_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12512__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11720__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12276__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ _02002_ _02450_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__nor2_1
XANTENNA__09141__A1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08480_ _03427_ _03428_ _03429_ _03430_ net692 net711 vssd1 vssd1 vccd1 vccd1 _03431_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06647__X _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12028__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11272__Y _05972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07431_ net760 _02381_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11713__B _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07362_ final_design.cpu.reg_window\[835\] final_design.cpu.reg_window\[867\] net944
+ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ final_design.CPU_instr_adr\[3\] _04023_ net1050 vssd1 vssd1 vccd1 vccd1 _00214_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11787__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07293_ final_design.cpu.reg_window\[5\] final_design.cpu.reg_window\[37\] net904
+ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09032_ _03960_ _03962_ net627 vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08514__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11539__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12200__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold300 final_design.cpu.reg_window\[701\] vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 final_design.cpu.reg_window\[684\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12036__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout203_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 final_design.cpu.reg_window\[696\] vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08955__A1 final_design.CPU_instr_adr\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07302__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold333 final_design.cpu.reg_window\[152\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1083 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold344 final_design.cpu.reg_window\[746\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13316__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold355 final_design.cpu.reg_window\[962\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 final_design.cpu.reg_window\[373\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 final_design.cpu.reg_window\[658\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net805 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_4
Xhold388 final_design.cpu.reg_window\[604\] vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ net472 _04732_ net483 vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__o21a_1
Xhold399 final_design.cpu.reg_window\[394\] vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout813 net814 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1112_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout824 net826 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__clkbuf_4
Xfanout835 net840 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_37_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09345__S net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout846 net848 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09904__B1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout857 net877 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_4
X_09865_ _04781_ _04783_ net498 vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__a21oi_1
Xhold1000 final_design.cpu.reg_window\[488\] vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 net869 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout572_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout193_X net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1011 final_design.cpu.reg_window\[811\] vssd1 vssd1 vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 net886 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07915__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1022 final_design.uart.working_data\[3\] vssd1 vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09380__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08816_ _03759_ _03761_ _03764_ _03766_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__a31o_1
Xhold1033 final_design.cpu.reg_window\[539\] vssd1 vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06813__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11607__C net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1044 final_design.cpu.reg_window\[297\] vssd1 vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ _03357_ net443 net439 _03356_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__o22a_1
Xhold1055 final_design.cpu.reg_window\[327\] vssd1 vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 final_design.cpu.reg_window\[32\] vssd1 vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ net673 _01598_ final_design.CPU_instr_adr\[7\] vssd1 vssd1 vccd1 vccd1 _03698_
+ sky130_fd_sc_hd__a21o_1
Xhold1077 final_design.cpu.reg_window\[293\] vssd1 vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12267__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12951__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 final_design.cpu.reg_window\[563\] vssd1 vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 final_design.cpu.reg_window\[302\] vssd1 vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout837_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08678_ _03617_ net603 vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_159_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14104__RESET_B net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09683__A2 _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07629_ final_design.cpu.reg_window\[476\] final_design.cpu.reg_window\[508\] net875
+ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__mux2_1
XANTENNA__11623__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_46_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10640_ net67 _05382_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09868__X _04787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11778__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10571_ _05291_ _05294_ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__or3_1
XFILLER_0_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12310_ net1876 net210 net365 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13290_ clknet_leaf_3_clk _00521_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[278\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12241_ net583 _06171_ net514 net374 net1506 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__a32o_1
XFILLER_0_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09738__A3 _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06452__B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_163_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__A2 _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ net2061 net219 net381 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11950__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ _02095_ net815 vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_55_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07564__A _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11054_ _05776_ _05777_ net1557 net1046 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06709__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11702__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ _04703_ _04885_ _04906_ _04923_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__and4_1
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06467__X _01418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11956_ net597 _06118_ _06158_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_28_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10907_ final_design.CPU_instr_adr\[22\] _03879_ net1071 vssd1 vssd1 vccd1 vccd1
+ _05637_ sky130_fd_sc_hd__mux2_1
XANTENNA__08882__B1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11887_ net242 net2102 net276 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09778__X _04697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10838_ _05549_ _05551_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__nand2_1
X_13626_ clknet_leaf_160_clk _00857_ net1105 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[614\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09426__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12430__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10769_ _05497_ _05503_ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__or3_1
X_13557_ clknet_leaf_40_clk _00788_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[545\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12508_ _06170_ net348 net327 net1961 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13488_ clknet_leaf_114_clk _00719_ net1211 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[476\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12439_ net1738 net245 net335 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07296__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11941__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14109_ clknet_leaf_83_clk _01306_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07980_ _01909_ net620 vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__nor2_1
XANTENNA__06789__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06931_ net549 _01881_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09362__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ _04567_ _04568_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__or2_1
X_06862_ _01809_ _01810_ _01811_ _01812_ net785 net793 vssd1 vssd1 vccd1 vccd1 _01813_
+ sky130_fd_sc_hd__mux4_1
X_08601_ net622 _03550_ _02423_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08570__C1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09581_ _03134_ _03582_ _04499_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__and3_1
X_06793_ final_design.cpu.reg_window\[854\] final_design.cpu.reg_window\[886\] net905
+ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__mux2_1
XANTENNA__09114__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ _02361_ net624 vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_26_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09665__A2 _04301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08463_ _03408_ _03413_ net722 vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__mux2_1
XANTENNA__11443__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08873__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07414_ final_design.cpu.reg_window\[321\] final_design.cpu.reg_window\[353\] net936
+ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__mux2_1
X_08394_ _03341_ _03342_ _03343_ _03344_ net685 net706 vssd1 vssd1 vccd1 vccd1 _03345_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_169_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09417__A2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07345_ _01484_ _02295_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08752__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout418_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09200__Y _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ net767 _02226_ net754 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_171_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09015_ net630 _03947_ _03946_ net256 vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout206_X net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08928__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 net102 vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09864__A _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13150__RESET_B net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 final_design.VGA_data_control.data_to_VGA\[16\] vssd1 vssd1 vccd1 vccd1 net1494
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold152 final_design.VGA_data_control.ready_data\[9\] vssd1 vssd1 vccd1 vccd1 net1505
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 final_design.VGA_data_control.ready_data\[15\] vssd1 vssd1 vccd1 vccd1 net1516
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout787_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 final_design.VGA_data_control.ready_data\[28\] vssd1 vssd1 vccd1 vccd1 net1527
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 net138 vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_2
Xhold196 final_design.cpu.reg_window\[717\] vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1115_X net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout621 _02513_ vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_4
Xfanout632 net633 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_4
X_09917_ net486 _04407_ _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__o21ai_1
Xfanout643 _06123_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout654 _05849_ vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_4
XANTENNA_fanout575_X net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout954_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout665 _05142_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_97_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout676 net678 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_4
Xfanout687 net689 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__buf_4
X_09848_ net735 _04763_ _04765_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__or3_2
XANTENNA__11160__A1 final_design.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout698 _01787_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_126_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ net75 _04186_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10432__A_N net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11810_ _06091_ net292 vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__nand2_1
XANTENNA__07323__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11999__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ net224 net2018 net416 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11672_ net230 net2307 net297 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10623_ net1017 _05365_ _05366_ net1042 net1377 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13411_ clknet_leaf_2_clk _00642_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[399\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10018__A3 _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08662__B _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_21_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13342_ clknet_leaf_146_clk _00573_ net1127 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[330\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input83_A memory_size[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10554_ net677 _05287_ _05300_ net979 _05299_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__o221a_1
XFILLER_0_64_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13273_ clknet_leaf_164_clk _00504_ net1085 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[261\]
+ sky130_fd_sc_hd__dfrtp_1
X_10485_ net90 final_design.VGA_adr\[0\] vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12224_ net592 _06152_ net519 net379 net1606 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__a32o_1
XANTENNA__07846__X _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11923__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09592__A1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__X _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ net188 net2451 net386 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__mux2_1
X_11106_ _05819_ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12086_ net586 _06039_ net515 net394 net1701 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__a32o_1
XANTENNA__10432__B _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_88_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11037_ net88 net1058 vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_34_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14026__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12988_ net1330 _00219_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06638__A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07202__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11939_ _06140_ net278 net408 net2381 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12651__B2 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13609_ clknet_leaf_84_clk _00840_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[597\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08572__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07130_ final_design.cpu.reg_window\[779\] final_design.cpu.reg_window\[811\] net938
+ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07061_ final_design.cpu.reg_window\[141\] final_design.cpu.reg_window\[173\] net913
+ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07269__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10717__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09583__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12314__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ final_design.cpu.reg_window\[209\] final_design.cpu.reg_window\[241\] net827
+ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_79_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06914_ final_design.cpu.reg_window\[210\] final_design.cpu.reg_window\[242\] net901
+ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09702_ _04092_ _04312_ _04298_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__o21ai_2
X_07894_ final_design.cpu.reg_window\[87\] final_design.cpu.reg_window\[119\] net843
+ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__mux2_1
XANTENNA__11142__A1 _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07346__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09886__A2 _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09633_ _04550_ _04551_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__xor2_1
X_06845_ net762 _01795_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout270_A net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout368_A net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09564_ _03132_ net442 net441 _03133_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__a2bb2o_1
X_06776_ final_design.cpu.reg_window\[278\] final_design.cpu.reg_window\[310\] net905
+ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08515_ final_design.cpu.reg_window\[130\] final_design.cpu.reg_window\[162\] net858
+ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__mux2_1
XANTENNA__13749__RESET_B net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09495_ _02607_ net445 net440 _02606_ _04413_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_121_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08310__A2 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08446_ final_design.cpu.reg_window\[68\] final_design.cpu.reg_window\[100\] net858
+ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08377_ _02240_ net610 vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout702_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07328_ final_design.cpu.reg_window\[132\] final_design.cpu.reg_window\[164\] net939
+ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08074__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07259_ _02204_ _02209_ net764 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12158__A0 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10270_ final_design.uart.BAUD_counter\[25\] final_design.uart.BAUD_counter\[24\]
+ _05128_ final_design.uart.BAUD_counter\[26\] vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__a31o_1
XFILLER_0_108_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10092__X _05008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout440 _04095_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_4
Xfanout451 _04069_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_4
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_2
X_13960_ clknet_leaf_119_clk _01191_ net1199 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[948\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout473 _03485_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_2
Xfanout484 net489 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12330__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout495 _03453_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_2
X_12911_ clknet_leaf_157_clk _00149_ net1112 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11684__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13891_ clknet_leaf_4_clk _01122_ net1096 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[879\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11364__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12842_ clknet_leaf_86_clk _00080_ net1249 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06458__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07053__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12633__B2 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07988__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11724_ net589 net423 _06220_ net297 net1566 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__a32o_1
XANTENNA__13419__RESET_B net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__A _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11655_ net189 net640 vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12397__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13072__RESET_B net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input86_X net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10606_ net98 final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__or2_1
X_11586_ net190 net644 vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10427__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13001__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10537_ _05283_ _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__nand2_1
X_13325_ clknet_leaf_139_clk _00556_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[313\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07812__B2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10468_ net677 _05216_ _05219_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__o21a_1
X_13256_ clknet_leaf_118_clk _00487_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[244\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12207_ net575 _06135_ net510 net376 net1777 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__a32o_1
XANTENNA__12134__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13187_ clknet_leaf_7_clk _00418_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[175\]
+ sky130_fd_sc_hd__dfrtp_1
X_10399_ net255 _05182_ net1048 net134 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07228__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12138_ net219 net2335 net385 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12069_ net583 _05911_ net514 net394 net1968 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_1_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07423__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07879__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06630_ _01577_ _01578_ _01579_ _01580_ net789 net806 vssd1 vssd1 vccd1 vccd1 _01581_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06551__A1 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13842__RESET_B net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06561_ final_design.cpu.reg_window\[285\] final_design.cpu.reg_window\[317\] net959
+ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__mux2_1
X_08300_ final_design.cpu.reg_window\[841\] final_design.cpu.reg_window\[873\] net843
+ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09280_ _02641_ _04172_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__xnor2_1
X_06492_ final_design.cpu.reg_window\[926\] final_design.cpu.reg_window\[958\] net931
+ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08231_ final_design.cpu.reg_window\[779\] final_design.cpu.reg_window\[811\] net857
+ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__mux2_1
XANTENNA__11721__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12309__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08162_ final_design.cpu.reg_window\[207\] final_design.cpu.reg_window\[239\] net824
+ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10938__A1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07113_ net750 net673 net671 _02061_ _01821_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_113_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08093_ final_design.cpu.reg_window\[460\] final_design.cpu.reg_window\[492\] net848
+ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload50 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_77_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07044_ net896 _01988_ _01994_ _01981_ _01982_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a32oi_1
Xclkload61 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_63_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload72 clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__inv_6
XANTENNA__08522__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload83 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_3_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload94 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 clkload94/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12044__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1025_A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12560__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08995_ final_design.CPU_instr_adr\[15\] _03791_ vssd1 vssd1 vccd1 vccd1 _03930_
+ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_10_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout485_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07946_ net618 _02894_ _02895_ net554 vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a211oi_1
XANTENNA__08758__A final_design.CPU_instr_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11666__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ _02824_ _02825_ _02826_ _02827_ net693 net702 vssd1 vssd1 vccd1 vccd1 _02828_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_162_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout652_A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout273_X net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07381__B _02330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07965__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09616_ _02867_ net441 vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__nand2_1
X_06828_ final_design.cpu.reg_window\[661\] final_design.cpu.reg_window\[693\] net965
+ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__mux2_1
XANTENNA__12615__A1 final_design.reqhand.data_from_UART\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_06759_ net760 _01709_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__or2_1
X_09547_ net483 _04377_ _04116_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout917_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__A0 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09478_ net468 _03639_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__or2_1
XANTENNA__07601__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11631__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08429_ final_design.cpu.reg_window\[581\] final_design.cpu.reg_window\[613\] net821
+ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ net1535 net178 net312 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__mux2_1
Xclkload0 clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_151_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10929__A1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ _04280_ _04285_ net660 vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10322_ net1729 net1022 net999 final_design.data_from_mem\[7\] vssd1 vssd1 vccd1
+ vccd1 _00079_ sky130_fd_sc_hd__a22o_1
X_13110_ clknet_leaf_130_clk _00341_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_14090_ clknet_leaf_71_clk _01287_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06741__A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08432__S net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13041_ clknet_leaf_91_clk _00272_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_10253_ net1724 _05119_ _05121_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12551__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input46_A mem_adr_start[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ final_design.uart.BAUD_counter\[1\] final_design.uart.BAUD_counter\[7\] final_design.uart.BAUD_counter\[6\]
+ final_design.uart.BAUD_counter\[0\] vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__or4b_1
Xfanout1202 net1209 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__buf_2
Xfanout1213 net1215 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__clkbuf_4
Xfanout1224 net1256 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__buf_2
Xfanout1235 net1238 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_4
Xfanout1246 net1256 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout270 net271 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_6
Xfanout281 net282 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_4
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_4
X_13943_ clknet_leaf_137_clk _01174_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[931\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13874_ clknet_leaf_26_clk _01105_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[862\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14178__Q final_design.VGA_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ net1367 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12606__B2 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09483__A0 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12756_ _06351_ _06385_ _06344_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06475__X _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12082__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11707_ net201 net634 vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__and2_1
X_12687_ final_design.VGA_data_control.ready_data\[31\] net1032 net987 final_design.data_from_mem\[31\]
+ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10438__A _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11638_ net437 net594 _06176_ net302 net1485 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__a32o_1
XFILLER_0_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11569_ net569 net420 _06140_ net303 net2108 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__a32o_1
XANTENNA__11593__A1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold707 final_design.cpu.reg_window\[77\] vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13308_ clknet_leaf_144_clk _00539_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[296\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold718 final_design.cpu.reg_window\[73\] vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 final_design.cpu.reg_window\[440\] vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09538__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13239_ clknet_leaf_144_clk _00470_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[227\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14041__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09962__A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07800_ net721 _02744_ net731 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__o21a_1
X_08780_ _03690_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10901__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07731_ final_design.cpu.reg_window\[218\] final_design.cpu.reg_window\[250\] net872
+ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__mux2_1
XANTENNA__11648__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07662_ final_design.cpu.reg_window\[286\] final_design.cpu.reg_window\[318\] net849
+ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06613_ _01560_ _01561_ _01562_ _01563_ net786 net794 vssd1 vssd1 vccd1 vccd1 _01564_
+ sky130_fd_sc_hd__mux4_1
X_09401_ net264 _04311_ _04313_ _04319_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__and4_1
XFILLER_0_149_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07593_ net626 _02540_ _02541_ _02502_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_172_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09332_ _04196_ _04250_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__and2_1
X_06544_ _01463_ _01474_ _01480_ _01482_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__or4_4
XANTENNA__09474__A0 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06826__A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12073__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08744__C _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09263_ net99 _04181_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__or2_2
XFILLER_0_145_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09202__A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06475_ final_design.data_from_mem\[18\] net981 _01425_ vssd1 vssd1 vccd1 vccd1 _01426_
+ sky130_fd_sc_hd__o21a_4
XANTENNA__12039__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06545__B net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08214_ _03164_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09194_ net603 _04111_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08145_ net890 _03095_ _03084_ _03083_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__09777__A1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout400_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1142_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08252__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ net606 _03022_ _02998_ net549 vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__o211a_1
XANTENNA__06686__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09529__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07027_ final_design.cpu.reg_window\[78\] final_design.cpu.reg_window\[110\] net926
+ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__mux2_1
XANTENNA__11336__A1 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1028_X net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_164_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout867_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 final_design.cpu.reg_window\[14\] vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 final_design.cpu.reg_window\[1\] vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 final_design.reqhand.instruction\[21\] vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ net627 _03912_ net256 vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__a21o_1
Xhold45 final_design.uart.working_data\[1\] vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 final_design.VGA_data_control.data_to_VGA\[10\] vssd1 vssd1 vccd1 vccd1 net1409
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07392__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 final_design.VGA_data_control.data_to_VGA\[31\] vssd1 vssd1 vccd1 vccd1 net1420
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 final_design.cpu.reg_window\[734\] vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _02876_ _02877_ _02878_ _02879_ net682 net704 vssd1 vssd1 vccd1 vccd1 _02880_
+ sky130_fd_sc_hd__mux4_1
Xhold89 final_design.VGA_data_control.data_to_VGA\[24\] vssd1 vssd1 vccd1 vccd1 net1442
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__C1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10940_ _05602_ _05622_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10871_ _05562_ _05578_ _05579_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__or3_1
XFILLER_0_151_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12610_ net1439 net1009 net995 final_design.data_from_mem\[28\] vssd1 vssd1 vccd1
+ vccd1 _01303_ sky130_fd_sc_hd__a22o_1
XANTENNA_input100_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12064__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13590_ clknet_leaf_124_clk _00821_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[578\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11272__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12541_ _06204_ net352 net323 net2183 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_6__f_clk_X clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12472_ _06254_ net502 net331 net2178 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14211_ net1280 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
X_11423_ net2060 net209 net311 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ clknet_leaf_75_clk _01316_ net1253 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11354_ _04381_ _04384_ net660 vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08162__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10705__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ final_design.VGA_data_control.h_count\[3\] net1061 _05158_ vssd1 vssd1 vccd1
+ vccd1 _05159_ sky130_fd_sc_hd__or3b_1
X_14073_ clknet_leaf_52_clk _01270_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11285_ final_design.data_from_mem\[16\] _02062_ _02509_ _05912_ _05917_ vssd1 vssd1
+ vccd1 vccd1 _05983_ sky130_fd_sc_hd__a41o_1
XFILLER_0_120_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11327__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12524__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10236_ final_design.uart.BAUD_counter\[13\] _05109_ net810 vssd1 vssd1 vccd1 vccd1
+ _05111_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09782__A _04697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13024_ clknet_leaf_36_clk _00255_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input49_X net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11878__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1010 _06295_ vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_2
Xfanout1021 _05170_ vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__buf_2
X_10167_ _05040_ _05057_ _05060_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[7\]
+ sky130_fd_sc_hd__and3_1
Xfanout1032 _06298_ vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_4
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__buf_4
Xfanout1054 _01371_ vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__buf_4
Xfanout1065 final_design.uart.receiving vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_2
Xfanout1076 net1080 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_4
X_10098_ net1062 _05012_ net1061 final_design.VGA_data_control.h_count\[3\] vssd1
+ vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__a211o_1
Xfanout1087 net1095 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__clkbuf_4
Xfanout1098 net1099 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10440__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07929__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13926_ clknet_leaf_168_clk _01157_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[914\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13434__RESET_B net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13857_ clknet_leaf_154_clk _01088_ net1116 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[845\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06601__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12808_ net1396 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13788_ clknet_leaf_153_clk _01019_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[776\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12739_ _05058_ _06366_ _06376_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__and3_1
XFILLER_0_155_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11802__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold504 final_design.cpu.reg_window\[941\] vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold515 final_design.cpu.reg_window\[996\] vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07865__S0 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold526 final_design.cpu.reg_window\[693\] vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold537 final_design.cpu.reg_window\[401\] vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold548 final_design.cpu.reg_window\[561\] vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ _04438_ _04112_ _04436_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__or3b_1
Xhold559 final_design.cpu.reg_window\[494\] vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11318__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12515__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08901_ _03665_ _03667_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_70_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11869__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ net475 _04797_ _04798_ net493 vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__a31o_1
XANTENNA__07617__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11286__X _05984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ net632 _02508_ net260 _03782_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a211o_1
XANTENNA__12322__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1204 net116 vssd1 vssd1 vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07942__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1215 final_design.cpu.reg_window\[308\] vssd1 vssd1 vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11446__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08763_ _02391_ _02393_ final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 _03714_
+ sky130_fd_sc_hd__a21boi_1
XANTENNA__10350__B net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08101__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout183_A _06067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09144__C1 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13175__RESET_B net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07714_ final_design.cpu.reg_window\[923\] final_design.cpu.reg_window\[955\] net882
+ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux2_1
X_08694_ _02772_ _03296_ _03593_ _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__and4_1
X_07645_ final_design.cpu.reg_window\[732\] final_design.cpu.reg_window\[764\] net874
+ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1092_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08755__B _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11462__A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07576_ net726 _02526_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07151__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10057__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06527_ _01379_ net1052 net1007 net1004 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__or4_1
X_09315_ _04232_ _04233_ net476 vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06458_ net1073 net1053 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__nand2_2
X_09246_ _04158_ _04164_ _04133_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09177_ _02544_ _04094_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1145_X net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08128_ final_design.cpu.reg_window\[13\] final_design.cpu.reg_window\[45\] net830
+ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08973__A2 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08059_ net717 _03003_ net730 vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12506__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ _05773_ _05776_ _05791_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__or3_1
XANTENNA__13945__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11908__Y _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ _04936_ _04937_ _04938_ net733 vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a211o_4
XANTENNA__10541__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06736__A1 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06831__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__A _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11972_ _06174_ net287 net405 net1660 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13711_ clknet_leaf_94_clk _00942_ net1226 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[699\]
+ sky130_fd_sc_hd__dfrtp_1
X_10923_ _05650_ _05651_ _05631_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11372__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06595__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13642_ clknet_leaf_1_clk _00873_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[630\]
+ sky130_fd_sc_hd__dfrtp_1
X_10854_ net78 _05548_ _05551_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12898__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10048__A1 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__B1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13573_ clknet_leaf_4_clk _00804_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[561\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10785_ net676 _05509_ _05518_ net974 _05520_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__o221a_1
XANTENNA__09453__A3 _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12524_ _06186_ net356 net329 net1656 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12455_ net1699 net193 net335 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07297__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11406_ net655 net176 vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12386_ net1742 net195 net270 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14125_ clknet_leaf_74_clk final_design.vga.v_next_count\[5\] net1252 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[5\] sky130_fd_sc_hd__dfrtp_4
X_11337_ _01722_ net649 _06028_ net652 net663 vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14056_ clknet_leaf_47_clk _00018_ net1148 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11268_ net667 _03932_ net739 vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ net1349 _00238_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[27\]
+ sky130_fd_sc_hd__dfrtp_2
X_10219_ final_design.uart.BAUD_counter\[6\] _05098_ _05100_ net811 vssd1 vssd1 vccd1
+ vccd1 _00034_ sky130_fd_sc_hd__o211a_1
XANTENNA__12142__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11199_ net667 _03992_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11720__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09677__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09141__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ clknet_leaf_25_clk _01140_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[897\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07688__C1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10597__S net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07430_ _02377_ _02378_ _02379_ _02380_ net781 net800 vssd1 vssd1 vccd1 vccd1 _02381_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_46_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11282__A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11713__C net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07361_ net764 _02305_ net756 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09100_ _04021_ _04022_ net260 vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07292_ final_design.cpu.reg_window\[69\] final_design.cpu.reg_window\[101\] net904
+ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08591__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09031_ _03731_ _03961_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10626__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12317__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08404__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold301 final_design.cpu.reg_window\[461\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09601__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold312 final_design.cpu.reg_window\[538\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 final_design.cpu.reg_window\[78\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 final_design.cpu.reg_window\[846\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__A2 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold345 final_design.cpu.reg_window\[471\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 final_design.cpu.reg_window\[155\] vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 final_design.cpu.reg_window\[765\] vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 final_design.cpu.reg_window\[526\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 final_design.cpu.reg_window\[854\] vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net477 _04795_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout803 net805 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_4
Xfanout814 _04039_ vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout825 net826 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout398_A net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout836 net840 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout847 net848 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12052__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09864_ _04112_ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__or2_1
Xfanout858 net860 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1105_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout869 net876 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_4
Xhold1001 final_design.cpu.reg_window\[311\] vssd1 vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 final_design.cpu.reg_window\[46\] vssd1 vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11176__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08815_ final_design.CPU_instr_adr\[22\] _01756_ _03755_ _03756_ vssd1 vssd1 vccd1
+ vccd1 _03766_ sky130_fd_sc_hd__a31o_1
XANTENNA__09380__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1023 final_design.cpu.reg_window\[552\] vssd1 vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 final_design.cpu.reg_window\[300\] vssd1 vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _04340_ _04709_ _04713_ _04348_ _04708_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__a32o_1
XANTENNA__06813__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1045 final_design.cpu.reg_window\[36\] vssd1 vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11891__S net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout186_X net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout565_A _05869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1056 final_design.cpu.reg_window\[808\] vssd1 vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 final_design.cpu.reg_window\[937\] vssd1 vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ final_design.CPU_instr_adr\[7\] net674 _01598_ vssd1 vssd1 vccd1 vccd1 _03697_
+ sky130_fd_sc_hd__and3_1
Xhold1078 final_design.reqhand.instruction\[5\] vssd1 vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 final_design.cpu.reg_window\[43\] vssd1 vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ net603 _03617_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_159_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1095_X net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07628_ final_design.cpu.reg_window\[284\] final_design.cpu.reg_window\[316\] net874
+ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__mux2_1
XANTENNA__12019__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12991__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07559_ _02094_ _02509_ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__or2_2
XFILLER_0_49_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10570_ _05314_ _05315_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__and2_1
XANTENNA__09840__B1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ _03638_ _04146_ _03637_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12240_ net576 _06170_ net510 net372 net1605 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout987_X net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12171_ net2329 net244 net382 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11122_ _01372_ _04993_ net1046 _05837_ net1354 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__o32a_1
Xhold890 final_design.cpu.reg_window\[624\] vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
X_11053_ _05757_ _05775_ _05172_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__a21o_1
XANTENNA__06709__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08254__S0 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ _04918_ _04921_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06895__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11955_ _06156_ net285 net409 net2283 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10906_ _05634_ _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08882__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11886_ net228 net2292 net274 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ clknet_leaf_167_clk _00856_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[613\]
+ sky130_fd_sc_hd__dfrtp_1
X_10837_ net78 _05548_ _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13556_ clknet_leaf_103_clk _00787_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[544\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08634__A1 _03296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10768_ _05496_ _05477_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__and2b_1
XANTENNA__12430__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09300__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12507_ _06169_ net351 net328 net1655 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12137__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10441__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__A _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13487_ clknet_leaf_91_clk _00718_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[475\]
+ sky130_fd_sc_hd__dfrtp_1
X_10699_ _05402_ _05421_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__or2_1
X_12438_ net1831 net238 net336 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12194__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12369_ net1786 net224 net270 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__mux2_1
XANTENNA__07296__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06930__Y _01881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14108_ clknet_leaf_83_clk _01305_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08350__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14039_ clknet_leaf_50_clk _00031_ net1155 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_06930_ net750 net673 net671 net761 _01821_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_38_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06861_ final_design.cpu.reg_window\[532\] final_design.cpu.reg_window\[564\] net948
+ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08600_ net622 _03550_ _02423_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__a21o_1
X_06792_ net767 _01742_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__nor2_1
X_09580_ _03164_ _04498_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11457__A0 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ _02361_ net612 vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08462_ _03409_ _03410_ _03411_ _03412_ net691 net702 vssd1 vssd1 vccd1 vccd1 _03413_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08873__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07413_ _02362_ _02363_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__or2_1
X_08393_ final_design.cpu.reg_window\[902\] final_design.cpu.reg_window\[934\] net831
+ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09417__A3 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07344_ final_design.data_from_mem\[11\] final_design.reqhand.instruction\[11\] net981
+ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08525__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12421__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08752__C _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07275_ _02222_ _02223_ _02224_ _02225_ net777 net792 vssd1 vssd1 vccd1 vccd1 _02226_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12047__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout313_A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06873__A_N _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09014_ _02448_ _03945_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08389__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11886__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold120 final_design.cpu.reg_window\[206\] vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 final_design.VGA_data_control.data_to_VGA\[12\] vssd1 vssd1 vccd1 vccd1 net1484
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1222_A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold142 _01331_ vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold153 final_design.cpu.reg_window\[715\] vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 final_design.VGA_data_control.data_to_VGA\[3\] vssd1 vssd1 vccd1 vccd1 net1517
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10291__S0 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold175 final_design.cpu.reg_window\[204\] vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 final_design.uart.BAUD_counter\[13\] vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 final_design.VGA_data_control.ready_data\[1\] vssd1 vssd1 vccd1 vccd1 net1550
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _05844_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_4
Xfanout611 net615 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09338__C1 _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout622 net624 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_4
X_09916_ net486 _04646_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__nand2_1
Xfanout633 _02506_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_2
Xfanout644 _06123_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_4
XANTENNA__12488__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout655 _05849_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_4
XANTENNA__10499__A1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout666 _03649_ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_4
Xfanout677 net678 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11696__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ _04763_ _04765_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout688 net690 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_4
XANTENNA_fanout947_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 net701 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ net737 _04681_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__and3_2
XANTENNA__07604__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08729_ final_design.CPU_instr_adr\[15\] _01967_ vssd1 vssd1 vccd1 vccd1 _03680_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ net240 net2531 net418 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11671_ net680 _05848_ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13410_ clknet_leaf_20_clk _00641_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[398\]
+ sky130_fd_sc_hd__dfrtp_1
X_10622_ _05347_ _05364_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09813__A0 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12412__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09120__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11620__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13341_ clknet_leaf_14_clk _00572_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[329\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10553_ net1067 _05295_ net1014 final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1
+ vccd1 _05300_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_8_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06722__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input76_A memory_size[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13272_ clknet_leaf_137_clk _00503_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[260\]
+ sky130_fd_sc_hd__dfrtp_1
X_10484_ _04880_ net253 _04990_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12176__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12223_ net589 _06151_ net516 net378 net1695 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__a32o_1
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13278__RESET_B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09592__A2 _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ net190 net2432 net386 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__mux2_1
XANTENNA__08170__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ net813 _05823_ _05825_ net976 vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08227__S0 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12085_ net571 _06032_ net506 net392 net2029 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__a32o_1
XANTENNA__12479__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11036_ _05722_ _05739_ _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11544__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12987_ net1329 _00218_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07107__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11938_ _06139_ net287 net409 net2428 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__a22o_1
XANTENNA__12651__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07202__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__B2 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11869_ _06109_ net290 net522 net2527 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13608_ clknet_leaf_126_clk _00839_ net1193 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[596\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12403__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07815__C1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13539_ clknet_leaf_7_clk _00770_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[527\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12094__C net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07060_ final_design.cpu.reg_window\[205\] final_design.cpu.reg_window\[237\] net913
+ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07269__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11719__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07962_ final_design.cpu.reg_window\[17\] final_design.cpu.reg_window\[49\] net827
+ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__mux2_1
X_09701_ net484 _04619_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__and2_1
X_06913_ final_design.cpu.reg_window\[18\] final_design.cpu.reg_window\[50\] net901
+ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11678__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07346__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07893_ _02840_ _02841_ _02842_ _02843_ net690 net710 vssd1 vssd1 vccd1 vccd1 _02844_
+ sky130_fd_sc_hd__mux4_1
X_09632_ net83 _04191_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_74_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06844_ _01791_ _01792_ _01793_ _01794_ net785 net803 vssd1 vssd1 vccd1 vccd1 _01795_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09563_ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__inv_2
XANTENNA__11454__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06775_ final_design.cpu.reg_window\[342\] final_design.cpu.reg_window\[374\] net905
+ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout263_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08514_ final_design.cpu.reg_window\[194\] final_design.cpu.reg_window\[226\] net858
+ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_162_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09494_ _02608_ _04087_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08445_ _03392_ _03393_ _03394_ _03395_ net691 net711 vssd1 vssd1 vccd1 vccd1 _03396_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11850__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout430_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10694__A1_N net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1172_A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08376_ _03324_ _03325_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__or2_2
X_07327_ final_design.cpu.reg_window\[196\] final_design.cpu.reg_window\[228\] net939
+ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__mux2_1
XANTENNA__10405__B2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08074__A2 _03022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06704__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07258_ _02205_ _02206_ _02207_ _02208_ net778 net793 vssd1 vssd1 vccd1 vccd1 _02209_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_30_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout897_A _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07189_ _02136_ _02137_ _02138_ _02139_ net780 net792 vssd1 vssd1 vccd1 vccd1 _02140_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08457__S0 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 net431 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_4
Xfanout441 _04094_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_4
Xfanout452 _04069_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout463 _03519_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_92_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout474 net475 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12330__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout485 net489 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__clkbuf_4
X_12910_ clknet_leaf_156_clk _00148_ net1114 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11645__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout496 net497 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
X_13890_ clknet_leaf_14_clk _01121_ net1103 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[878\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07334__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ clknet_leaf_72_clk _00079_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11364__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07196__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11723_ net187 net636 vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__and2_1
XANTENNA__11841__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06943__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09121__Y _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11654_ net586 net423 _06184_ net301 net1718 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12397__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10605_ net98 final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11585_ net429 net578 _06148_ net304 net1956 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__a32o_1
XFILLER_0_88_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09785__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13324_ clknet_leaf_121_clk _00555_ net1197 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[312\]
+ sky130_fd_sc_hd__dfrtp_1
X_10536_ net62 _05282_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13255_ clknet_leaf_8_clk _00486_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[243\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10467_ net813 _05217_ _05218_ net975 vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__o22a_1
XANTENNA__10724__A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12206_ net577 _06134_ net512 net377 net1649 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__a32o_1
XANTENNA__09565__A2 _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13186_ clknet_leaf_29_clk _00417_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[174\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10398_ _03549_ _05181_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__or2_1
X_12137_ net244 net2393 net386 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12068_ net573 _05905_ net509 net392 net1706 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__a32o_1
X_11019_ _01359_ _03837_ net1072 vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__mux2_1
XANTENNA__12150__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06649__A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10332__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07423__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07244__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12085__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06560_ final_design.cpu.reg_window\[349\] final_design.cpu.reg_window\[381\] net959
+ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09312__X _04231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06491_ final_design.cpu.reg_window\[990\] final_design.cpu.reg_window\[1022\] net930
+ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ final_design.cpu.reg_window\[843\] final_design.cpu.reg_window\[875\] net857
+ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08161_ final_design.cpu.reg_window\[15\] final_design.cpu.reg_window\[47\] net824
+ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__mux2_1
XANTENNA__10399__B1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09695__A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07112_ net750 net673 _01851_ _02061_ _01821_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__o221a_1
XFILLER_0_160_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08092_ final_design.cpu.reg_window\[268\] final_design.cpu.reg_window\[300\] net846
+ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload40 clknet_leaf_146_clk vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__clkinv_4
X_07043_ net769 _01993_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload51 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_42_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12325__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload62 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__inv_6
Xclkload73 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_77_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload84 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload95 clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 clkload95/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11899__A0 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11363__A2 _05143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09961__C1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08994_ _03925_ _03929_ final_design.CPU_instr_adr\[16\] net1026 vssd1 vssd1 vccd1
+ vccd1 _00227_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_103_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07945_ net608 _02894_ _02869_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout380_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__A1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08758__B _02330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__A3 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09206__Y _04125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07876_ final_design.cpu.reg_window\[532\] final_design.cpu.reg_window\[564\] net867
+ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07154__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ net498 _04533_ _04231_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__o21ba_1
X_06827_ final_design.cpu.reg_window\[725\] final_design.cpu.reg_window\[757\] net964
+ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout266_X net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout645_A _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09546_ net492 _04368_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__and2_1
XANTENNA__12076__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06993__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06758_ _01705_ _01706_ _01707_ _01708_ net778 net798 vssd1 vssd1 vccd1 vccd1 _01709_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11823__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ net533 _02325_ net532 net531 net460 net468 vssd1 vssd1 vccd1 vccd1 _04396_
+ sky130_fd_sc_hd__mux4_1
X_06689_ final_design.cpu.reg_window\[217\] final_design.cpu.reg_window\[249\] net952
+ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12091__A3 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08428_ final_design.cpu.reg_window\[645\] final_design.cpu.reg_window\[677\] net821
+ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12379__A1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload1 clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__inv_6
X_08359_ final_design.cpu.reg_window\[839\] final_design.cpu.reg_window\[871\] net856
+ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11370_ net664 _06055_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10321_ net1499 net1022 net999 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1
+ vccd1 _00078_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10544__A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11339__C1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13040_ clknet_leaf_108_clk _00271_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10252_ final_design.uart.BAUD_counter\[19\] _05119_ net809 vssd1 vssd1 vccd1 vccd1
+ _05121_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12000__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ final_design.uart.BAUD_counter\[3\] final_design.uart.BAUD_counter\[2\] final_design.uart.BAUD_counter\[5\]
+ final_design.uart.BAUD_counter\[4\] vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__or4b_1
Xfanout1203 net1209 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__clkbuf_4
Xfanout1214 net1215 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__clkbuf_4
Xfanout1225 net1239 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__clkbuf_4
Xfanout1236 net1238 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input39_A mem_adr_start[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1247 net1248 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__clkbuf_4
Xfanout260 net261 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout271 net273 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_31_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12303__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_4
X_13942_ clknet_leaf_125_clk _01173_ net1191 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[930\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07064__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13873_ clknet_leaf_109_clk _01104_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[861\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07999__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12067__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12824_ net1375 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10617__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11814__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12755_ _06344_ _06351_ _06385_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__and3_1
XANTENNA__10617__B2 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09483__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06916__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11706_ net426 net571 _06211_ net295 net1957 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12686_ _06330_ net1458 net993 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10438__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11637_ net221 net641 vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14210__1279 vssd1 vssd1 vccd1 vccd1 _14210__1279/HI net1279 sky130_fd_sc_hd__conb_1
XFILLER_0_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11568_ net205 net642 vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07341__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13307_ clknet_leaf_136_clk _00538_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[295\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold708 final_design.cpu.reg_window\[648\] vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11593__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10519_ _05249_ _05264_ _05263_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__a21oi_1
Xhold719 final_design.cpu.reg_window\[770\] vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12145__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10454__A _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11499_ net816 _05842_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_139_Left_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07239__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13238_ clknet_leaf_130_clk _00469_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[226\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09538__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11345__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09962__B _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ clknet_leaf_107_clk _00400_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[157\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10553__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10901__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07730_ final_design.cpu.reg_window\[26\] final_design.cpu.reg_window\[58\] net870
+ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07661_ final_design.cpu.reg_window\[350\] final_design.cpu.reg_window\[382\] net849
+ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_148_Left_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09400_ net499 _04298_ _04301_ _04074_ _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__o221a_1
X_06612_ final_design.cpu.reg_window\[540\] final_design.cpu.reg_window\[572\] net951
+ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07592_ net612 _02540_ _02515_ _02502_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09331_ net89 _04195_ net91 vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11291__Y _05989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06543_ _01474_ _01482_ _01481_ _01464_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_48_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11805__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09474__A1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10629__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09262_ net98 _04180_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__and2_1
X_06474_ final_design.reqhand.instruction\[18\] net984 vssd1 vssd1 vccd1 vccd1 _01425_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_118_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10348__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06545__C _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08213_ _03162_ _03163_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_138_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09193_ _03617_ net666 vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__or2_4
X_12785__16 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__inv_2
XFILLER_0_62_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout226_A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11033__A1 _05673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12230__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08144_ _03089_ _03094_ net727 vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_157_Left_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload140 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 clkload140/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_116_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12055__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ net550 _03024_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_31_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1135_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07026_ final_design.cpu.reg_window\[142\] final_design.cpu.reg_window\[174\] net926
+ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11894__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout595_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_164_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold13 final_design.cpu.reg_window\[24\] vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 net131 vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09591__C _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08977_ _02456_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout762_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 net149 vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 final_design.VGA_data_control.data_to_VGA\[8\] vssd1 vssd1 vccd1 vccd1 net1399
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 final_design.VGA_data_control.data_to_VGA\[23\] vssd1 vssd1 vccd1 vccd1 net1410
+ sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ final_design.cpu.reg_window\[150\] final_design.cpu.reg_window\[182\] net819
+ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__mux2_1
XANTENNA__09388__S1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold68 final_design.reqhand.instruction\[25\] vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 final_design.VGA_data_control.data_to_VGA\[1\] vssd1 vssd1 vccd1 vccd1 net1432
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09162__B1 _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_166_Left_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07859_ _02806_ _02807_ _02808_ _02809_ net693 net712 vssd1 vssd1 vccd1 vccd1 _02810_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10870_ _05600_ _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09529_ net496 _04439_ _04447_ _04231_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ _06203_ net351 net324 net1933 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12471_ _06131_ net344 net331 net2152 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14210_ net1279 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XFILLER_0_136_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11422_ net1691 net211 net312 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__mux2_1
XANTENNA__12221__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06752__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11575__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14141_ clknet_leaf_75_clk _01315_ net1245 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11353_ _01660_ net650 _06042_ net653 net664 vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10304_ final_design.VGA_data_control.data_to_VGA\[31\] final_design.VGA_data_control.data_to_VGA\[30\]
+ final_design.VGA_data_control.data_to_VGA\[29\] final_design.VGA_data_control.data_to_VGA\[28\]
+ net1063 net1062 vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__mux4_1
X_14072_ clknet_leaf_52_clk _01269_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11284_ _03613_ _05913_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13023_ clknet_leaf_133_clk _00254_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10235_ _05109_ _05110_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__nor2_1
Xfanout1000 _05167_ vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__buf_2
Xfanout1011 _06295_ vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__buf_2
XANTENNA__09127__X _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1022 net1023 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__buf_2
X_10166_ _05054_ _05058_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__nand2_1
Xfanout1033 _06298_ vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_2
Xfanout1044 _04994_ vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__buf_4
Xfanout1055 net1056 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__buf_2
Xfanout1066 net1069 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__buf_2
XANTENNA__12288__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1077 net1080 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_2
X_10097_ net1063 net1062 vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__and2_1
Xfanout1088 net1095 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__clkbuf_2
Xfanout1099 net1104 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_2
XFILLER_0_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ clknet_leaf_149_clk _01156_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[913\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload4_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13856_ clknet_leaf_38_clk _01087_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[844\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06486__X _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12807_ net1407 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09303__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13474__RESET_B net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13787_ clknet_leaf_155_clk _01018_ net1115 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[775\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10999_ _04042_ _05715_ _05724_ _04040_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12738_ net967 _06377_ _06378_ net808 net2567 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__a32o_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12669_ final_design.VGA_data_control.ready_data\[22\] net1032 net987 final_design.data_from_mem\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12212__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold505 final_design.cpu.reg_window\[789\] vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 final_design.cpu.reg_window\[581\] vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07865__S1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold527 final_design.cpu.reg_window\[799\] vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 final_design.cpu.reg_window\[659\] vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 final_design.cpu.reg_window\[281\] vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
X_08900_ final_design.CPU_instr_adr\[26\] net1029 _03842_ _03845_ vssd1 vssd1 vccd1
+ vccd1 _00237_ sky130_fd_sc_hd__a22o_1
X_09880_ net477 _04795_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_70_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07617__S1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08831_ net632 _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__nor2_1
XANTENNA__11727__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1205 final_design.cpu.reg_window\[411\] vssd1 vssd1 vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 final_design.VGA_adr\[0\] vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07942__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08762_ net1031 _02361_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12279__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09144__B1 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07713_ final_design.cpu.reg_window\[987\] final_design.cpu.reg_window\[1019\] net881
+ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08693_ _03359_ _03425_ _03636_ _03643_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__and4_1
XFILLER_0_170_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12294__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout176_A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07644_ net722 _02594_ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11462__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07575_ _02522_ _02523_ _02524_ _02525_ net688 net709 vssd1 vssd1 vccd1 vccd1 _02526_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout343_A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1085_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09314_ net540 net539 net538 net537 net457 net466 vssd1 vssd1 vccd1 vccd1 _04233_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__10057__A2 _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06526_ _01465_ _01468_ _01475_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__or3_2
XANTENNA__11254__A1 _02030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11889__S net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09245_ _04132_ _04162_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06457_ wb_manage.BUSY_O net1073 net34 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout510_A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08670__A2 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout229_X net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout608_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12203__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08263__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ _03631_ _03650_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11557__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08127_ final_design.cpu.reg_window\[77\] final_design.cpu.reg_window\[109\] net830
+ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1040_X net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09883__A _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08058_ net725 _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__nor2_1
XANTENNA__12580__Y _06295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout977_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ final_design.cpu.reg_window\[719\] final_design.cpu.reg_window\[751\] net907
+ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__mux2_1
XANTENNA__09907__C1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10822__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A0 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ _04936_ _04937_ _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11637__B net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ _06173_ net281 net404 net1654 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__a22o_1
XANTENNA__12285__A3 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13710_ clknet_leaf_116_clk _00941_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[698\]
+ sky130_fd_sc_hd__dfrtp_1
X_10922_ net83 net1060 vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07342__S net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06595__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13641_ clknet_leaf_85_clk _00872_ net1235 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[629\]
+ sky130_fd_sc_hd__dfrtp_1
X_10853_ final_design.CPU_instr_adr\[20\] _03893_ net1070 vssd1 vssd1 vccd1 vccd1
+ _05585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11245__B2 _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ clknet_leaf_98_clk _00803_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[560\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09989__A2 _04773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10784_ net974 _05519_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12523_ _06185_ net353 net329 net2001 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12454_ net1928 net195 net335 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__mux2_1
XANTENNA__08173__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08949__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11405_ net599 _06087_ _06088_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__and3_2
XFILLER_0_22_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12385_ net1798 _06017_ net273 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14124_ clknet_leaf_74_clk final_design.vga.v_next_count\[4\] net1252 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11336_ final_design.data_from_mem\[23\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06028_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_91_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14055_ clknet_leaf_47_clk _00016_ net1148 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11267_ final_design.data_from_mem\[15\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1
+ _05967_ sky130_fd_sc_hd__a21o_2
XFILLER_0_24_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10508__B1 final_design.CPU_instr_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13006_ net1348 _00237_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_10218_ _05099_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11198_ final_design.data_from_mem\[7\] final_design.reqhand.data_from_UART\[7\]
+ net253 vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__mux2_2
XANTENNA__08202__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11181__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ final_design.VGA_data_control.h_count\[0\] _05013_ vssd1 vssd1 vccd1 vccd1
+ _05048_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12276__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908_ clknet_leaf_102_clk _01139_ net1188 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[896\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09141__A3 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12681__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08348__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07252__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13839_ clknet_leaf_90_clk _01070_ net1233 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[827\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07360_ net771 _02310_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08637__C1 _01938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11787__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07291_ _02239_ _02240_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_135_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11502__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09030_ _03688_ _03689_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10626__B final_design.VGA_adr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold302 final_design.cpu.reg_window\[969\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08404__A2 _03352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12200__A3 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold313 final_design.cpu.reg_window\[234\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 net159 vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 final_design.cpu.reg_window\[861\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 final_design.cpu.reg_window\[919\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 final_design.cpu.reg_window\[1022\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11297__X _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09932_ _04179_ _04850_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__or2_1
Xhold368 final_design.cpu.reg_window\[476\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold379 final_design.cpu.reg_window\[605\] vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout804 net805 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__buf_2
Xfanout815 _02392_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09365__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout826 net829 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout837 net840 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_2
X_09863_ _04690_ _04779_ net484 vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__mux2_1
Xfanout848 net855 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_2
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net860 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_4
X_08814_ _03764_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__inv_2
Xhold1002 final_design.cpu.reg_window\[315\] vssd1 vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 final_design.cpu.reg_window\[817\] vssd1 vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1024 final_design.cpu.reg_window\[120\] vssd1 vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ net483 _04712_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__nand2_1
XANTENNA__09380__A3 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1035 final_design.cpu.reg_window\[106\] vssd1 vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 final_design.cpu.reg_window\[954\] vssd1 vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ final_design.CPU_instr_adr\[8\] _02186_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__and2_1
Xhold1057 final_design.cpu.reg_window\[619\] vssd1 vssd1 vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1068 final_design.cpu.reg_window\[822\] vssd1 vssd1 vccd1 vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout460_A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 final_design.cpu.reg_window\[632\] vssd1 vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12267__A3 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09668__B2 _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_X net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08676_ _03625_ _03626_ _03619_ _03621_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__o211a_2
XANTENNA__08258__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11192__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07627_ final_design.cpu.reg_window\[348\] final_design.cpu.reg_window\[380\] net874
+ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout725_A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07558_ _01998_ _02028_ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__nor2_1
XANTENNA__12424__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11778__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06509_ net1053 net1006 net1003 _01376_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_3_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07489_ _02185_ _02186_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08643__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1255_X net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11412__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09228_ _03638_ _04146_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09159_ net623 _03550_ _01597_ _02423_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14113__RESET_B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12170_ net2030 net237 net380 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__mux2_1
X_11121_ _01373_ net1045 _04993_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10552__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold880 final_design.cpu.reg_window\[928\] vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 final_design.cpu.reg_window\[571\] vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07337__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ _05757_ _05775_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__nor2_1
XANTENNA__08254__S1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06709__A2 _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ _04919_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nand2_1
XANTENNA__11702__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09405__X _04324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__A3 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954_ _06155_ net286 net409 net2124 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__a22o_1
XANTENNA__08168__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07072__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10905_ _05629_ _05633_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__and2b_1
XFILLER_0_157_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ net230 net2379 net276 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__mux2_1
XANTENNA_output108_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_103_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11218__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13624_ clknet_leaf_131_clk _00855_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[612\]
+ sky130_fd_sc_hd__dfrtp_1
X_10836_ _05567_ _05568_ _05548_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12415__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13555_ clknet_leaf_34_clk _00786_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[543\]
+ sky130_fd_sc_hd__dfrtp_1
X_10767_ _05479_ _05498_ _05478_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__and3b_1
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10286__X _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10727__A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11322__S net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12430__A3 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12506_ _06168_ net347 net327 net1726 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__a22o_1
XANTENNA__06645__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10441__A2 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__B _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13486_ clknet_leaf_114_clk _00717_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[474\]
+ sky130_fd_sc_hd__dfrtp_1
X_10698_ _05436_ _05437_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10446__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12437_ net1828 net223 net335 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09595__B1 _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12368_ net1838 net240 net272 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14107_ clknet_leaf_71_clk _01304_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_112_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11319_ net743 _03886_ _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11941__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11558__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12153__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10462__A _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ net2072 _05875_ net366 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14038_ clknet_leaf_51_clk _00028_ net1155 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_06860_ final_design.cpu.reg_window\[596\] final_design.cpu.reg_window\[628\] net948
+ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__mux2_1
X_06791_ _01738_ _01739_ _01740_ _01741_ net774 net795 vssd1 vssd1 vccd1 vccd1 _01742_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12249__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08530_ _03468_ _03469_ _03480_ net891 vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08461_ final_design.cpu.reg_window\[516\] final_design.cpu.reg_window\[548\] net860
+ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11209__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07412_ net532 _02361_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__and2_1
XFILLER_0_174_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12406__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08392_ final_design.cpu.reg_window\[966\] final_design.cpu.reg_window\[998\] net830
+ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07343_ _02281_ _02282_ _02293_ net899 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_73_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12328__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07274_ final_design.cpu.reg_window\[6\] final_design.cpu.reg_window\[38\] net914
+ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09013_ net630 _03944_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_171_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08389__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1048_A _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12185__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 final_design.cpu.reg_window\[556\] vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 net130 vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08541__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold132 final_design.cpu.reg_window\[208\] vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 final_design.reqhand.instruction\[27\] vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 final_design.VGA_data_control.data_to_VGA\[21\] vssd1 vssd1 vccd1 vccd1 net1507
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11468__A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11932__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold165 final_design.cpu.reg_window\[205\] vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 net106 vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10291__S1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold187 final_design.cpu.reg_window\[196\] vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09338__B1 _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout601 _05199_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__buf_6
Xhold198 final_design.cpu.reg_window\[713\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 net615 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_2
X_09915_ net537 net536 net534 net533 net454 net463 vssd1 vssd1 vccd1 vccd1 _04834_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout623 net624 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__buf_1
XANTENNA__11145__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout634 net635 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_4
XANTENNA_fanout296_X net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 _06123_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_2
Xfanout656 net658 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__buf_4
Xfanout667 _02512_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_4
XANTENNA__11696__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ _04673_ _04764_ net448 vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13506__RESET_B net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout678 _04989_ vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__buf_2
Xfanout689 net690 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__buf_2
X_09777_ _04046_ _04350_ _04682_ _04695_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_126_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06989_ net547 _01939_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout842_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _01363_ _01968_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__nor2_1
XANTENNA__09510__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11999__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08659_ net262 _03596_ _03609_ _03595_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_1_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08864__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11670_ net817 _02358_ net815 vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__nand3_1
XFILLER_0_138_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10621_ _05347_ _05364_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09401__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__A1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10959__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13340_ clknet_leaf_147_clk _00571_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[328\]
+ sky130_fd_sc_hd__dfrtp_1
X_10552_ net978 _05298_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__nand2_1
XANTENNA__11620__A1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06722__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13271_ clknet_leaf_142_clk _00502_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[259\]
+ sky130_fd_sc_hd__dfrtp_1
X_10483_ net36 _05220_ _05228_ _05229_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12222_ net584 _06150_ net514 net378 net2003 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__a32o_1
XANTENNA_input69_A memory_size[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11923__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ net192 net2495 net384 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__mux2_1
XANTENNA__09592__A3 _04508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11104_ net972 _05822_ _05824_ net970 vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__o22a_1
XANTENNA__07067__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12084_ net2406 net392 net500 _06025_ vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__a22o_1
XANTENNA__08227__S1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11035_ _05720_ _05739_ _05738_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_34_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10895__C1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11439__A1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12986_ net1328 _00217_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11937_ _06138_ net281 net408 net2238 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_165_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_165_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11868_ net426 net200 net563 net520 net1983 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__a32o_1
XANTENNA__07530__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10819_ _05551_ _05552_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11560__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13607_ clknet_leaf_10_clk _00838_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[595\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12148__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11799_ net654 net565 net195 vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__and3_1
XANTENNA__09804__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13538_ clknet_leaf_23_clk _00769_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[526\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07910__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13469_ clknet_leaf_12_clk _00700_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[457\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10904__B _05629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11375__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07961_ final_design.cpu.reg_window\[81\] final_design.cpu.reg_window\[113\] net828
+ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__mux2_1
XANTENNA__11127__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09700_ _04457_ _04618_ net472 vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__mux2_1
X_06912_ final_design.cpu.reg_window\[82\] final_design.cpu.reg_window\[114\] net901
+ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__mux2_1
XANTENNA__11678__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ final_design.cpu.reg_window\[407\] final_design.cpu.reg_window\[439\] net852
+ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08597__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07346__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09631_ net737 _04546_ _04549_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__and3_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06843_ final_design.cpu.reg_window\[404\] final_design.cpu.reg_window\[436\] net953
+ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__mux2_1
XANTENNA_wire529_X net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ _04186_ _04480_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_104_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06774_ _01718_ _01722_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_104_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09205__B _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08513_ final_design.cpu.reg_window\[2\] final_design.cpu.reg_window\[34\] net865
+ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10102__A1 final_design.VGA_data_control.v_count\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_172_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ _04208_ _04210_ net468 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_156_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_156_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout256_A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08444_ final_design.cpu.reg_window\[388\] final_design.cpu.reg_window\[420\] net859
+ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06845__A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08059__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08375_ _03297_ _03322_ net537 vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__a21o_1
XANTENNA__12058__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout423_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1165_A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07326_ final_design.cpu.reg_window\[4\] final_design.cpu.reg_window\[36\] net939
+ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__mux2_1
XANTENNA__10405__A2 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06704__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11897__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07257_ final_design.cpu.reg_window\[519\] final_design.cpu.reg_window\[551\] net937
+ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout211_X net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07188_ final_design.cpu.reg_window\[9\] final_design.cpu.reg_window\[41\] net924
+ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__mux2_1
XANTENNA__11366__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_A _01419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__S1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1218_X net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10614__A2_N net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 net421 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_4
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout431 _05847_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11926__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout442 net445 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_4
Xfanout453 net454 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_4
Xfanout464 net465 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_2
Xfanout475 _03485_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12330__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07615__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout486 net489 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09731__B1 _04648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ net735 _04744_ _04747_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__o21a_1
XANTENNA__11645__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout497 _03419_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_4
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10341__B2 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ clknet_leaf_72_clk _00078_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_147_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_147_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11722_ net435 net591 _06219_ net297 net2236 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07196__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08446__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07350__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06943__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11653_ net190 net640 vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__and2_1
X_10604_ net254 _04787_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__and2b_1
XANTENNA__12397__A2 _06268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ net192 net643 vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13323_ clknet_leaf_20_clk _00554_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[311\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10535_ net62 _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13254_ clknet_leaf_171_clk _00485_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[242\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10466_ net68 net971 net969 final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1
+ _05218_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10724__B _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11357__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12205_ net575 _06133_ net510 net377 net1817 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__a32o_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13185_ clknet_leaf_159_clk _00416_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[173\]
+ sky130_fd_sc_hd__dfrtp_1
X_10397_ _03648_ _05180_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__or2_4
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12136_ net237 net2454 net384 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__mux2_1
XANTENNA__09970__B1 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11109__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__C1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ net573 _05898_ net508 net393 net1816 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_53_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09722__A0 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ final_design.CPU_instr_adr\[27\] net1014 _05742_ net1067 vssd1 vssd1 vccd1
+ vccd1 _05743_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07959__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13010__RESET_B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08210__A _02000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10332__B2 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12085__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_138_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_138_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12969_ clknet_leaf_46_clk _00207_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.uart.bits_received\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06490_ final_design.cpu.reg_window\[798\] final_design.cpu.reg_window\[830\] net931
+ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08160_ final_design.cpu.reg_window\[79\] final_design.cpu.reg_window\[111\] net824
+ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10399__B2 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07111_ final_design.reqhand.instruction\[12\] net986 _02060_ vssd1 vssd1 vccd1 vccd1
+ _02062_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09695__B _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08091_ final_design.cpu.reg_window\[332\] final_design.cpu.reg_window\[364\] net846
+ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__mux2_1
XANTENNA__06698__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11510__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload30 clknet_leaf_157_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__clkinv_4
Xclkload41 clknet_leaf_148_clk vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__clkinv_4
X_07042_ _01989_ _01990_ _01991_ _01992_ net781 net801 vssd1 vssd1 vccd1 vccd1 _01993_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08091__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13851__RESET_B net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06604__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload52 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload63 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__clkinv_8
Xclkload74 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 clkload74/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07016__A1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload85 clknet_leaf_136_clk vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__inv_6
XANTENNA__12903__Q net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload96 clknet_leaf_145_clk vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__inv_6
XANTENNA__13169__RESET_B net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12560__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ net257 _03927_ net1026 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_166_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07944_ _01755_ net608 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07875_ final_design.cpu.reg_window\[596\] final_design.cpu.reg_window\[628\] net866
+ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10323__B2 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout373_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06826_ net765 _01776_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__or2_1
X_09614_ net494 _04491_ _04227_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ _02936_ net446 net442 _02932_ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_129_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06757_ final_design.cpu.reg_window\[919\] final_design.cpu.reg_window\[951\] net918
+ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout540_A _02126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09476_ _04393_ _04394_ net479 vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__mux2_1
X_06688_ final_design.cpu.reg_window\[25\] final_design.cpu.reg_window\[57\] net952
+ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__mux2_1
XANTENNA__09492__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08427_ final_design.cpu.reg_window\[709\] final_design.cpu.reg_window\[741\] net821
+ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10097__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1070_X net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout805_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1168_X net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08358_ net718 _03302_ net730 vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__o21a_1
XFILLER_0_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload2 clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__inv_6
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11587__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07309_ final_design.cpu.reg_window\[581\] final_design.cpu.reg_window\[613\] net904
+ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08452__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08289_ final_design.cpu.reg_window\[9\] final_design.cpu.reg_window\[41\] net842
+ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__mux2_1
XANTENNA__10825__A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11420__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10320_ net1542 net1025 net1002 final_design.data_from_mem\[5\] vssd1 vssd1 vccd1
+ vccd1 _00077_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10251_ _05119_ _05120_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12551__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ _05069_ _05071_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout962_X net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1204 net1209 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1215 net1216 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1226 net1239 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__clkbuf_2
Xfanout1237 net1238 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__clkbuf_4
Xfanout250 _04986_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_4
Xfanout1248 net1255 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__clkbuf_4
Xfanout261 _03654_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_6
X_13941_ clknet_leaf_25_clk _01172_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[929\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout283 _06228_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_4
Xfanout294 _06228_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06613__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13872_ clknet_leaf_111_clk _01103_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[860\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07191__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12067__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ net1360 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08684__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12754_ _06344_ _06351_ _06384_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__or3_1
XANTENNA__06485__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09483__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06916__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11705_ net203 net634 vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__and2_1
X_12685_ final_design.VGA_data_control.ready_data\[30\] net1034 net989 final_design.data_from_mem\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__a22o_1
XANTENNA__11290__A2 _05984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input91_X net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11636_ net426 net569 _06175_ net299 net1582 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__a32o_1
XFILLER_0_170_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11567_ net578 net422 _06139_ net304 net2056 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06932__B _01881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ net1479 net1045 net1017 _05266_ vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07341__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13306_ clknet_leaf_163_clk _00537_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[294\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08994__B2 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold709 final_design.cpu.reg_window\[380\] vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11498_ net681 _06116_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__nand2_1
XANTENNA__10454__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13237_ clknet_leaf_40_clk _00468_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[225\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09538__A3 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10449_ net1491 net1048 _05208_ net248 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_161_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09943__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13168_ clknet_leaf_105_clk _00399_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[156\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11750__A0 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10553__B2 final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ net1751 net190 net390 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12161__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ clknet_leaf_13_clk _00330_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07108__X _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ _01507_ net613 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_140_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06611_ final_design.cpu.reg_window\[604\] final_design.cpu.reg_window\[636\] net951
+ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07591_ net612 _02540_ _02515_ _02503_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__o211a_1
X_09330_ net733 _04248_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__or2_2
XANTENNA__11505__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06542_ _01463_ _01474_ _01482_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__or3_4
XFILLER_0_133_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10629__B final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09474__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09261_ net96 net97 _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06473_ final_design.cpu.reg_window\[286\] final_design.cpu.reg_window\[318\] net930
+ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08212_ net604 _03160_ _03135_ net545 vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09192_ _03617_ net666 vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__nor2_2
XFILLER_0_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11569__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08143_ _03090_ _03091_ _03092_ _03093_ net685 net706 vssd1 vssd1 vccd1 vccd1 _03094_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout219_A _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08074_ net617 _03022_ _03023_ net550 vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__a211oi_2
Xclkload130 clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 clkload130/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload141 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 clkload141/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__08115__A _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07025_ final_design.cpu.reg_window\[206\] final_design.cpu.reg_window\[238\] net926
+ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_168_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_129_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1030_A _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1128_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12533__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout490_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout588_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 final_design.cpu.reg_window\[23\] vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09591__D _04508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08976_ _01911_ _01912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__and2b_1
Xhold25 net171 vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12985__RESET_B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07165__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold36 net144 vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 final_design.VGA_data_control.data_to_VGA\[9\] vssd1 vssd1 vccd1 vccd1 net1400
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 final_design.reqhand.instruction\[22\] vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ final_design.cpu.reg_window\[214\] final_design.cpu.reg_window\[246\] net819
+ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__mux2_1
XANTENNA__12297__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold69 net123 vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout755_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08596__S0 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ final_design.cpu.reg_window\[404\] final_design.cpu.reg_window\[436\] net872
+ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06809_ final_design.cpu.reg_window\[213\] final_design.cpu.reg_window\[245\] net963
+ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__mux2_1
X_07789_ final_design.cpu.reg_window\[345\] final_design.cpu.reg_window\[377\] net863
+ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout922_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09528_ _04436_ _04446_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ _04107_ _04377_ _04376_ net483 vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_137_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09870__C1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12470_ _06130_ net344 net331 net2038 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11421_ net2201 net213 net313 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12221__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14140_ clknet_leaf_76_clk net1257 net1253 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.h_count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11352_ final_design.data_from_mem\[25\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06042_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10303_ final_design.VGA_data_control.h_count\[3\] _05156_ final_design.VGA_data_control.h_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10783__B2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11980__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14071_ clknet_leaf_52_clk _01268_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11283_ net437 net593 _05981_ net318 net1662 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__a32o_1
XANTENNA__12770__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ clknet_leaf_21_clk _00253_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input51_A mem_adr_start[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ final_design.uart.BAUD_counter\[12\] _05108_ net810 vssd1 vssd1 vccd1 vccd1
+ _05110_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12524__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07087__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06739__B1 _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1001 _05167_ vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__buf_2
Xfanout1012 _06295_ vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_2
X_10165_ _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__inv_2
Xfanout1023 _05166_ vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__buf_2
Xfanout1034 _06298_ vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1045 net1047 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__buf_2
Xfanout1056 net1057 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_1
XANTENNA__12288__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ final_design.VGA_data_control.h_count\[0\] net1063 vssd1 vssd1 vccd1 vccd1
+ _05012_ sky130_fd_sc_hd__or2_1
Xfanout1067 net1069 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__clkbuf_4
Xfanout1078 net1080 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__clkbuf_4
Xfanout1089 net1095 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13924_ clknet_leaf_106_clk _01155_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[912\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06767__X _01718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13855_ clknet_leaf_135_clk _01086_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[843\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12806_ net1404 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11552__C net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10998_ _05722_ _05723_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__or2_1
X_13786_ clknet_leaf_162_clk _01017_ net1105 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[774\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09456__A2 _04302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12737_ _05058_ _06373_ _06376_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__a21o_1
XANTENNA__08664__B1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__A2 _05960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10471__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12668_ _06321_ net1507 net991 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11619_ net245 net638 vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__and2_1
XANTENNA__12156__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12599_ net1390 net1010 net996 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1
+ vccd1 _01292_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07110__Y _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08511__S0 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold506 final_design.cpu.reg_window\[980\] vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11971__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold517 final_design.cpu.reg_window\[543\] vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 final_design.cpu.reg_window\[82\] vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold539 final_design.cpu.reg_window\[421\] vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12515__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08830_ _03779_ _03780_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06825__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1206 wb_manage.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08761_ _01367_ _02361_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1217 final_design.cpu.reg_window\[407\] vssd1 vssd1 vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08578__S0 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07712_ final_design.cpu.reg_window\[795\] final_design.cpu.reg_window\[827\] net882
+ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__mux2_1
X_08692_ _03456_ _03457_ _03554_ _03639_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__and4_1
XFILLER_0_174_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06677__X _01628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07643_ _02590_ _02591_ _02592_ _02593_ net694 net713 vssd1 vssd1 vccd1 vccd1 _02594_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06902__B1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07574_ final_design.cpu.reg_window\[159\] final_design.cpu.reg_window\[191\] net841
+ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__mux2_1
XANTENNA__10905__A_N _05629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09313_ net545 net544 net543 net541 net458 net467 vssd1 vssd1 vccd1 vccd1 _04232_
+ sky130_fd_sc_hd__mux4_1
X_06525_ _01465_ _01468_ _01475_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__nor3_1
XANTENNA__11254__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12451__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout336_A _06282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09244_ _04162_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1078_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06456_ _01405_ _01406_ _01407_ _01396_ vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_118_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12203__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ _03631_ _03650_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout503_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1245_A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08126_ _03073_ _03074_ _03075_ _03076_ net685 net700 vssd1 vssd1 vccd1 vccd1 _03077_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11962__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ _03004_ _03005_ _03006_ _03007_ net682 net704 vssd1 vssd1 vccd1 vccd1 _03008_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12506__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07008_ _01955_ _01956_ _01957_ _01958_ net775 net796 vssd1 vssd1 vccd1 vccd1 _01959_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11918__B _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09383__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09458__A_N _04308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ _02459_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11970_ _06172_ net285 net405 net1561 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_16_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10921_ net83 net1060 vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__and2_1
XANTENNA__11653__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07241__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10852_ _04954_ net251 vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__nor2_1
X_13640_ clknet_leaf_127_clk _00871_ net1193 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[628\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10783_ final_design.CPU_instr_adr\[16\] net1013 _05516_ net1054 vssd1 vssd1 vccd1
+ vccd1 _05519_ sky130_fd_sc_hd__o22ai_1
X_13571_ clknet_leaf_7_clk _00802_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[559\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12765__A final_design.VGA_adr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _06184_ net356 net329 net1704 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input99_A memory_size[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12453_ net2149 net196 net338 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11404_ _04127_ _04176_ net664 vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12384_ net1790 net198 net272 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10300__S0 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11953__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14123_ clknet_leaf_74_clk final_design.vga.v_next_count\[3\] net1252 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[3\] sky130_fd_sc_hd__dfrtp_4
X_11335_ net745 _03869_ _06026_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14054_ clknet_leaf_47_clk _00015_ net1148 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06702__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11266_ net2365 net316 _05966_ net429 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10217_ final_design.uart.BAUD_counter\[6\] _05098_ vssd1 vssd1 vccd1 vccd1 _05099_
+ sky130_fd_sc_hd__and2_1
X_13005_ net1347 _00236_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[25\]
+ sky130_fd_sc_hd__dfrtp_2
X_11197_ net427 net573 _05905_ net315 net2130 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11181__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ _05012_ _05046_ _05047_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[1\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_27_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10079_ net1 _04995_ _04993_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_89_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07533__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ clknet_leaf_27_clk _01138_ net1139 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[895\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13832__Q final_design.cpu.reg_window\[820\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13838_ clknet_leaf_120_clk _01069_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[826\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12433__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13769_ clknet_leaf_84_clk _01000_ net1235 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[757\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_42_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07290_ _02239_ _02240_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10995__A1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09601__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11944__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 final_design.cpu.reg_window\[986\] vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold314 final_design.cpu.reg_window\[53\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 final_design.cpu.reg_window\[990\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 final_design.cpu.reg_window\[768\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 final_design.cpu.reg_window\[923\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 final_design.cpu.reg_window\[236\] vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ net95 _04178_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__nor2_1
XANTENNA_wire559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_3__f_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xhold369 final_design.cpu.reg_window\[157\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout805 net807 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_2
Xfanout816 _02295_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_4_7__f_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout827 net829 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_4
X_09862_ net487 _04683_ _04780_ _04055_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__a211o_1
Xfanout838 net839 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_4
Xfanout849 net851 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07915__A2 _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ final_design.CPU_instr_adr\[20\] _01823_ _03760_ vssd1 vssd1 vccd1 vccd1
+ _03764_ sky130_fd_sc_hd__a21bo_1
Xhold1003 final_design.cpu.reg_window\[367\] vssd1 vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09770__D1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1014 final_design.reqhand.instruction\[10\] vssd1 vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ _04710_ _04711_ net477 vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1025 final_design.cpu.reg_window\[96\] vssd1 vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 final_design.cpu.reg_window\[1020\] vssd1 vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1047 final_design.cpu.reg_window\[694\] vssd1 vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ final_design.CPU_instr_adr\[9\] net673 _01537_ vssd1 vssd1 vccd1 vccd1 _03695_
+ sky130_fd_sc_hd__and3_1
Xhold1058 final_design.cpu.reg_window\[920\] vssd1 vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07128__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08539__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1069 final_design.cpu.reg_window\[829\] vssd1 vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08675_ _02061_ _03616_ _01487_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10683__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07015__Y _01966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ _01570_ net613 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_159_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07557_ _02477_ _02505_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout620_A _02513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_X net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_33_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06508_ net1051 net1007 net1004 final_design.reqhand.instruction\[4\] vssd1 vssd1
+ vccd1 vccd1 _01459_ sky130_fd_sc_hd__o31a_1
XFILLER_0_124_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10435__B1 _05201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07488_ _02214_ _02437_ _02213_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a21oi_2
XANTENNA__06583__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06439_ wb_manage.BUSY_O net34 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__and2b_1
X_09227_ _03488_ _04145_ _03486_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09158_ _04075_ _04076_ net479 vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__mux2_1
XANTENNA__09053__B1 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06870__X _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10738__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10738__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11935__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08109_ final_design.cpu.reg_window\[652\] final_design.cpu.reg_window\[684\] net847
+ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09089_ _02300_ _02433_ _04012_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_114_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11120_ _05831_ _05835_ _05836_ _05830_ net2539 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__a32o_1
XANTENNA__07618__S net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold870 final_design.cpu.reg_window\[783\] vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 final_design.cpu.reg_window\[531\] vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ _05773_ _05774_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__or2_1
Xhold892 final_design.cpu.reg_window\[274\] vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
X_10002_ _04192_ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__and2_1
XANTENNA__12360__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08449__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07353__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11953_ _06154_ net293 net411 net2099 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12663__B2 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10904_ _05633_ _05629_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_28_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ _05848_ _06246_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_84_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13623_ clknet_leaf_136_clk _00854_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[611\]
+ sky130_fd_sc_hd__dfrtp_1
X_10835_ net78 net1055 vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_172_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09292__A0 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13554_ clknet_leaf_42_clk _00785_ net1150 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[542\]
+ sky130_fd_sc_hd__dfrtp_1
X_10766_ _05439_ _05501_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_41_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ _06167_ net348 net328 net1804 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10697_ net39 _05435_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__nor2_1
X_13485_ clknet_leaf_139_clk _00716_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[473\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12436_ net1861 net240 net337 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12434__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ net1627 net227 net272 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14106_ clknet_leaf_83_clk _01303_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07528__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11318_ net669 _03882_ net743 vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11558__B net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12298_ net2110 net228 net365 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10462__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14037_ clknet_leaf_51_clk _00017_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11249_ net655 net211 vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__and2_1
XANTENNA__12351__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08570__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06790_ final_design.cpu.reg_window\[662\] final_design.cpu.reg_window\[694\] net902
+ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__mux2_1
X_14244__1309 vssd1 vssd1 vccd1 vccd1 _14244__1309/HI net1309 sky130_fd_sc_hd__conb_1
XANTENNA__08359__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06668__A net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_11__f_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_106_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10665__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08460_ final_design.cpu.reg_window\[580\] final_design.cpu.reg_window\[612\] net858
+ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07411_ net532 _02361_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08391_ final_design.cpu.reg_window\[774\] final_design.cpu.reg_window\[806\] net835
+ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_102_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11513__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07342_ _02287_ _02292_ net762 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__mux2_1
XANTENNA__08094__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07273_ final_design.cpu.reg_window\[70\] final_design.cpu.reg_window\[102\] net914
+ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _02032_ _02033_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold100 final_design.reqhand.instruction\[15\] vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 final_design.cpu.reg_window\[202\] vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 final_design.VGA_data_control.ready_data\[29\] vssd1 vssd1 vccd1 vccd1 net1475
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold133 final_design.VGA_data_control.data_to_VGA\[6\] vssd1 vssd1 vccd1 vccd1 net1486
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11393__A1 final_design.data_from_mem\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold144 final_design.VGA_data_control.data_to_VGA\[26\] vssd1 vssd1 vccd1 vccd1 net1497
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold155 final_design.VGA_data_control.ready_data\[3\] vssd1 vssd1 vccd1 vccd1 net1508
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11468__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold166 final_design.cpu.reg_window\[991\] vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 final_design.reqhand.instruction\[7\] vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold188 final_design.uart.BAUD_counter\[28\] vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout602 _05199_ vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_2
X_09914_ _03422_ net444 net440 _03421_ _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__o221a_1
Xhold199 final_design.cpu.reg_window\[63\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout613 net615 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_2
XANTENNA__11145__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1110_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout624 net625 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout635 _06192_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12342__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1208_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 net648 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_6
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout657 net658 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__buf_2
XANTENNA__08010__B2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _03229_ _04503_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__or2_1
Xfanout668 _02512_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11696__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout570_A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 net680 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08269__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ _04409_ _04694_ _04689_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_126_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06988_ net750 net673 net671 net781 _01821_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__o221a_4
XTAP_TAPCELL_ROW_126_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _01939_ final_design.CPU_instr_adr\[16\] vssd1 vssd1 vccd1 vccd1 _03678_
+ sky130_fd_sc_hd__and2b_1
XANTENNA__12645__B2 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10656__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09889__A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _02642_ _03607_ _03608_ _02545_ _03604_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_166_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07901__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07609_ final_design.cpu.reg_window\[541\] final_design.cpu.reg_window\[573\] net878
+ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08589_ final_design.cpu.reg_window\[896\] final_design.cpu.reg_window\[928\] net862
+ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11423__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10620_ _05362_ _05363_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09813__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ _04042_ _05296_ _05297_ _05295_ net973 vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__a32o_1
XANTENNA__11620__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10482_ _05231_ _05232_ net1502 net1045 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_161_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09026__B1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13270_ clknet_leaf_128_clk _00501_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[258\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12221_ net586 _06149_ net515 net378 net1675 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__a32o_1
XANTENNA__11384__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ net194 net2309 net384 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__mux2_1
XANTENNA__10773__A_N net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08033__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ final_design.CPU_instr_adr\[31\] _03804_ net1072 vssd1 vssd1 vccd1 vccd1
+ _05824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09329__A1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12083_ net595 _06018_ net519 net395 net1908 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12333__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ _04421_ net252 vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__nor2_1
XANTENNA__07872__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07083__S net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12985_ net1327 _00216_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11936_ _06137_ net285 net409 net2316 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__a22o_1
XANTENNA__07811__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11867_ _06108_ net278 net520 net2273 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__a22o_1
X_13606_ clknet_leaf_170_clk _00837_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[594\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10818_ _05530_ _05533_ _05550_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_60_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11798_ net2491 net415 net292 _06018_ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13537_ clknet_leaf_157_clk _00768_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[525\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10749_ net74 net1056 vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07910__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13468_ clknet_leaf_147_clk _00699_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[456\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12419_ _06017_ net647 net359 _06280_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12164__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11375__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13399_ clknet_leaf_145_clk _00630_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[387\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14004__RESET_B net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07960_ net717 _02910_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__nor2_1
XANTENNA__11127__A1 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_4_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06911_ net758 _01861_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__nor2_1
XANTENNA__11678__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07891_ final_design.cpu.reg_window\[471\] final_design.cpu.reg_window\[503\] net852
+ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11508__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ _02868_ _04547_ _04548_ net448 vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__a211o_1
X_06842_ final_design.cpu.reg_window\[468\] final_design.cpu.reg_window\[500\] net949
+ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06554__A1 final_design.data_from_mem\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09561_ net73 _04185_ net74 vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__o21ai_1
X_06773_ _01723_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12627__B2 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08512_ final_design.cpu.reg_window\[66\] final_design.cpu.reg_window\[98\] net865
+ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09492_ net556 net555 net554 net553 net461 _03518_ vssd1 vssd1 vccd1 vccd1 _04411_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_19_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08443_ final_design.cpu.reg_window\[452\] final_design.cpu.reg_window\[484\] net859
+ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__mux2_1
XANTENNA__10648__A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11850__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout249_A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08059__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ net619 _03321_ _03323_ _02211_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12939__RESET_B net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07325_ final_design.cpu.reg_window\[68\] final_design.cpu.reg_window\[100\] net939
+ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__mux2_1
XANTENNA__11063__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout416_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1158_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ final_design.cpu.reg_window\[583\] final_design.cpu.reg_window\[615\] net915
+ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09559__A1 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07187_ final_design.cpu.reg_window\[73\] final_design.cpu.reg_window\[105\] net924
+ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout204_X net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11366__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07665__S0 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout410 net411 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_8
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_4
Xfanout432 net436 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_4
Xfanout443 net445 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_2
Xfanout454 net456 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout952_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11418__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 _03519_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_2
Xfanout476 net479 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08534__A2 _03481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09828_ _04182_ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12330__A3 _06268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout487 net489 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_2
Xfanout498 net499 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09759_ _04659_ _04677_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13380__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12770_ net1060 net808 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09495__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11721_ net188 net636 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__and2_1
XANTENNA__11661__B net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11652_ net429 net578 _06183_ net300 net2235 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__a32o_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10603_ _05329_ _05345_ _05344_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_80_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11583_ net425 net567 _06147_ net303 net2160 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__a32o_1
XANTENNA_input81_A memory_size[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13322_ clknet_leaf_4_clk _00553_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[310\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10534_ net677 _05269_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14243__1308 vssd1 vssd1 vccd1 vccd1 _14243__1308/HI net1308 sky130_fd_sc_hd__conb_1
XFILLER_0_162_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11389__A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10465_ final_design.CPU_instr_adr\[0\] net68 net1067 vssd1 vssd1 vccd1 vccd1 _05217_
+ sky130_fd_sc_hd__mux2_1
X_13253_ clknet_leaf_17_clk _00484_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[241\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11357__A1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10724__C net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12554__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12204_ _06132_ net502 net378 net2360 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10396_ _01481_ net734 net677 _05174_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__or4_2
X_13184_ clknet_leaf_37_clk _00415_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[172\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12135_ net223 net2295 net384 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__mux2_1
XANTENNA__09970__B2 _04066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12066_ net588 _05891_ net515 net394 net1884 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_53_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09722__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09183__C1 _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _05740_ _05741_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07959__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10332__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12609__B2 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12968_ clknet_leaf_52_clk _00206_ net1150 vssd1 vssd1 vccd1 vccd1 final_design.uart.bits_received\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07541__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11293__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ net179 _06248_ _06251_ net275 net2571 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__a32o_1
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12159__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12899_ clknet_leaf_68_clk _00137_ net1221 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07113__Y _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07110_ final_design.reqhand.instruction\[12\] net986 _02060_ vssd1 vssd1 vccd1 vccd1
+ _02061_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_43_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08090_ _02064_ net606 vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__nand2_1
XANTENNA__06681__A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06698__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload20 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__inv_6
X_07041_ final_design.cpu.reg_window\[654\] final_design.cpu.reg_window\[686\] net926
+ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload31 clknet_leaf_158_clk vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload42 clknet_leaf_150_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__clkinv_2
Xclkload53 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__bufinv_16
Xclkload64 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_77_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12545__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload75 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__09992__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload86 clknet_leaf_138_clk vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__inv_8
Xclkload97 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_149_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09961__A1 _04871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ _03927_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_166_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07943_ net888 _02875_ _02881_ _02887_ _02893_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__o32a_4
XTAP_TAPCELL_ROW_166_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout199_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13138__RESET_B net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ final_design.cpu.reg_window\[660\] final_design.cpu.reg_window\[692\] net866
+ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11520__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09613_ _04510_ _04511_ _04531_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07017__A _01967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06825_ _01772_ _01773_ _01774_ _01775_ net789 net806 vssd1 vssd1 vccd1 vccd1 _01776_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout366_A net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09477__A0 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ _02933_ net441 vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06756_ final_design.cpu.reg_window\[983\] final_design.cpu.reg_window\[1015\] net918
+ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12076__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07451__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06687_ final_design.cpu.reg_window\[89\] final_design.cpu.reg_window\[121\] net952
+ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__mux2_1
X_09475_ net538 net537 net536 net534 net457 net466 vssd1 vssd1 vccd1 vccd1 _04394_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout533_A _02294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09492__A3 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08426_ _03373_ _03374_ _03375_ _03376_ net684 net704 vssd1 vssd1 vccd1 vccd1 _03377_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10097__B net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08357_ net725 _03307_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout700_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1063_X net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11587__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07308_ _02255_ _02256_ _02257_ _02258_ net776 net795 vssd1 vssd1 vccd1 vccd1 _02259_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08452__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08288_ final_design.cpu.reg_window\[73\] final_design.cpu.reg_window\[105\] net842
+ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07239_ final_design.cpu.reg_window\[71\] final_design.cpu.reg_window\[103\] net916
+ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__mux2_1
XANTENNA__13979__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12536__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ net2561 _05118_ net809 vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12000__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13908__RESET_B net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _05067_ _05068_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__or3_1
XFILLER_0_121_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06766__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1205 net1209 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09407__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1216 net1217 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__clkbuf_2
Xfanout1227 net1239 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1238 net1239 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__clkbuf_2
Xfanout240 _05890_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout955_X net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout251 net255 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_4
Xfanout1249 net1251 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout273 _06278_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_8
X_13940_ clknet_leaf_101_clk _01171_ net1188 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[928\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout284 net287 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_4
Xfanout295 net298 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07810__S0 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06613__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ clknet_leaf_90_clk _01102_ net1233 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[859\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07191__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12822_ net1371 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11275__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12753_ _06351_ _06384_ _06344_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10288__A _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09483__A3 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11704_ net437 net594 _06210_ net298 net1846 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__a32o_1
XFILLER_0_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12684_ _06329_ net1403 net991 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11027__B1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11635_ net205 net638 vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input84_X net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08192__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07877__S0 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11566_ net207 net643 vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__and2_1
X_13305_ clknet_leaf_163_clk _00536_ net1085 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[293\]
+ sky130_fd_sc_hd__dfrtp_1
X_10517_ _05249_ _05265_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11497_ _02359_ _05838_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__nor2_1
XANTENNA__12527__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13236_ clknet_leaf_142_clk _00467_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[224\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10448_ net529 net602 vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_94_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13649__RESET_B net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12442__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ clknet_leaf_95_clk _00398_ net1226 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[155\]
+ sky130_fd_sc_hd__dfrtp_1
X_10379_ net22 net1037 net1020 net2572 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12118_ net2125 net192 net388 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11566__B net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13098_ clknet_leaf_0_clk _00329_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12049_ net2091 net194 net396 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06610_ final_design.cpu.reg_window\[668\] final_design.cpu.reg_window\[700\] net956
+ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__mux2_1
X_07590_ _02504_ net626 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__nor2_1
XANTENNA__08367__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06541_ _01482_ _01464_ _01473_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__and3b_1
XFILLER_0_133_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11805__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09474__A3 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09260_ net95 _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__and2_1
X_06472_ final_design.cpu.reg_window\[350\] final_design.cpu.reg_window\[382\] net930
+ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08211_ net616 _03160_ _03161_ net545 vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_172_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06693__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09191_ net481 _04083_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11521__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08142_ final_design.cpu.reg_window\[909\] final_design.cpu.reg_window\[941\] net832
+ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload120 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload120/Y sky130_fd_sc_hd__inv_8
XFILLER_0_114_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08073_ net606 _03022_ _02998_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_116_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload131 clknet_leaf_90_clk vssd1 vssd1 vccd1 vccd1 clkload131/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload142 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 clkload142/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__12518__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07024_ _01971_ _01972_ _01973_ _01974_ net781 net801 vssd1 vssd1 vccd1 vccd1 _01975_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_168_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07954__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1023_A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07446__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _03748_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout483_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 final_design.cpu.reg_window\[29\] vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 net120 vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 final_design.reqhand.instruction\[17\] vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ final_design.cpu.reg_window\[22\] final_design.cpu.reg_window\[54\] net819
+ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__mux2_1
Xhold48 final_design.reqhand.data_from_UART\[2\] vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 final_design.reqhand.instruction\[26\] vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08596__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ final_design.cpu.reg_window\[468\] final_design.cpu.reg_window\[500\] net868
+ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout271_X net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_A _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14242__1307 vssd1 vssd1 vccd1 vccd1 _14242__1307/HI net1307 sky130_fd_sc_hd__conb_1
XFILLER_0_39_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06808_ _01757_ _01758_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__nand2_1
X_07788_ _01660_ net611 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__nand2_1
XANTENNA__12954__RESET_B net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07181__S net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09527_ net474 _04336_ _04223_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__a21boi_2
X_06739_ net751 net674 _01504_ _01689_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout915_A net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09458_ _04308_ net473 _04054_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__and3b_1
XFILLER_0_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08409_ _02267_ net621 vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ net468 _03553_ _04061_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__or3_2
XFILLER_0_108_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11431__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11420_ net1801 net216 net312 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07859__S0 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09622__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11351_ net748 _03853_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06987__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10783__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12509__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10302_ final_design.VGA_data_control.data_to_VGA\[15\] final_design.VGA_data_control.data_to_VGA\[14\]
+ final_design.VGA_data_control.data_to_VGA\[13\] final_design.VGA_data_control.data_to_VGA\[12\]
+ net1063 net1062 vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__mux4_1
X_14070_ clknet_leaf_52_clk _01267_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.uart.working_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_89_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11282_ net658 net221 vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__and2_1
XANTENNA__12770__B net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13021_ clknet_leaf_11_clk _00252_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10233_ final_design.uart.BAUD_counter\[12\] _05108_ vssd1 vssd1 vccd1 vccd1 _05109_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07087__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__C1 _05901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07356__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input44_A mem_adr_start[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ final_design.VGA_data_control.VGA_request_address\[1\] final_design.VGA_data_control.VGA_request_address\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__and2_2
Xfanout1002 _05167_ vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09137__A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1013 net1014 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__buf_2
XANTENNA__08041__A _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1024 _05166_ vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1035 _06298_ vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1046 net1047 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_4
X_10095_ final_design.VGA_data_control.h_count\[5\] _05010_ vssd1 vssd1 vccd1 vccd1
+ _05011_ sky130_fd_sc_hd__or2_1
Xfanout1057 final_design.VGA_adr\[10\] vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__clkbuf_2
Xfanout1068 net1069 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__clkbuf_2
Xfanout1079 net1080 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_2
XANTENNA__07880__A _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13923_ clknet_leaf_6_clk _01154_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[911\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08900__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13854_ clknet_leaf_148_clk _01085_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[842\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_98_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08187__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ net1362 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ clknet_leaf_160_clk _01016_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[773\]
+ sky130_fd_sc_hd__dfrtp_1
X_10997_ _05717_ _05721_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_48_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07879__X _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12736_ _05059_ _06372_ _06376_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__or3b_1
XFILLER_0_84_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09861__B1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10471__A1 net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12667_ final_design.VGA_data_control.ready_data\[21\] net1032 net987 final_design.data_from_mem\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__a22o_1
XANTENNA__12437__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11618_ net573 net421 _06166_ net300 net1563 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__a32o_1
XFILLER_0_128_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12598_ net1384 net1009 net995 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1
+ vccd1 _01291_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08511__S1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07624__C1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11549_ net568 net420 _06130_ net303 net1796 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__a32o_1
XFILLER_0_41_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold507 final_design.cpu.reg_window\[957\] vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold518 final_design.cpu.reg_window\[703\] vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 final_design.cpu.reg_window\[674\] vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12790__21 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__inv_2
XFILLER_0_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ clknet_leaf_6_clk _00450_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[207\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12172__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199_ net1268 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XANTENNA__13412__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06825__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1207 final_design.VGA_data_control.state\[1\] vssd1 vssd1 vccd1 vccd1 net2560
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ _03709_ _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__and2b_1
Xhold1218 final_design.cpu.reg_window\[414\] vssd1 vssd1 vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11487__A0 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07711_ final_design.cpu.reg_window\[859\] final_design.cpu.reg_window\[891\] net882
+ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XANTENNA__08578__S1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08691_ _03554_ _03639_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__nand2_1
XANTENNA__11516__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07642_ final_design.cpu.reg_window\[924\] final_design.cpu.reg_window\[956\] net874
+ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08097__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06902__A1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07573_ final_design.cpu.reg_window\[223\] final_design.cpu.reg_window\[255\] net841
+ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__mux2_1
X_09312_ _04092_ _04218_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__or2_4
X_06524_ _01454_ _01455_ _01471_ _01472_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09243_ _04134_ _04159_ _04161_ _02995_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__a211o_1
X_06455_ _01405_ _01406_ _01407_ _01396_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout231_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout329_A net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09174_ net530 _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__nor2_1
XANTENNA__07030__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ final_design.cpu.reg_window\[269\] final_design.cpu.reg_window\[301\] net834
+ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1140_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10094__C _05008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1238_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08056_ final_design.cpu.reg_window\[146\] final_design.cpu.reg_window\[178\] net818
+ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07007_ final_design.cpu.reg_window\[911\] final_design.cpu.reg_window\[943\] net907
+ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__mux2_1
XANTENNA__09907__A1 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08266__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_X net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ _01855_ _01856_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__nand2b_1
XANTENNA__07904__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ final_design.cpu.reg_window\[535\] final_design.cpu.reg_window\[567\] net828
+ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08889_ net632 _03833_ _03834_ _03835_ net259 vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__a311o_1
XFILLER_0_99_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11426__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ _04550_ net247 net678 vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_168_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10150__B1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07241__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10851_ net1015 _05582_ _05583_ net1041 net1424 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__a32o_1
XFILLER_0_116_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout918_X net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_160_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13570_ clknet_leaf_28_clk _00801_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[558\]
+ sky130_fd_sc_hd__dfrtp_1
X_10782_ net972 _05516_ _05517_ net968 vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__o22a_1
XANTENNA__09843__B1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12765__B net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12521_ _06183_ net346 net327 net1579 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11650__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10453__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10566__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13994__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12452_ net2119 net198 net337 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11403_ net664 _06084_ _06086_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12383_ net1872 net200 net271 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__mux2_1
XANTENNA__10300__S1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14122_ clknet_leaf_74_clk final_design.vga.v_next_count\[2\] net1252 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[2\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_10_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11334_ net669 _03864_ net745 vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07621__A2 _02570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11397__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ clknet_leaf_48_clk _00014_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ net655 net582 net208 vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__and3_1
XANTENNA__10508__A2 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07086__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ net1346 _00235_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_10216_ _05098_ net812 _05097_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__and3b_1
X_11196_ net654 net237 vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__and2_1
XANTENNA__11181__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10147_ final_design.VGA_data_control.h_count\[0\] net1063 vssd1 vssd1 vccd1 vccd1
+ _05047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10078_ wb_manage.curr_state\[2\] wb_manage.curr_state\[1\] vssd1 vssd1 vccd1 vccd1
+ _04995_ sky130_fd_sc_hd__or2_1
XANTENNA__12130__A1 _06094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13906_ clknet_leaf_26_clk _01137_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[894\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07688__A2 _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12681__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07115__A _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10692__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13837_ clknet_leaf_127_clk _01068_ net1193 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[825\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10692__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_128_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13768_ clknet_leaf_118_clk _00999_ net1195 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[756\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08637__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09834__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09330__A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06648__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ _06355_ _06358_ _06356_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12167__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__10476__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13699_ clknet_leaf_1_clk _00930_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[687\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_135_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13664__RESET_B net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09062__A1 _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09476__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold304 final_design.cpu.reg_window\[594\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09329__X _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14241__1306 vssd1 vssd1 vccd1 vccd1 _14241__1306/HI net1306 sky130_fd_sc_hd__conb_1
Xhold315 final_design.cpu.reg_window\[1005\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08380__S net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold326 final_design.cpu.reg_window\[666\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 final_design.cpu.reg_window\[230\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 final_design.cpu.reg_window\[568\] vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ _04178_ _04829_ _04847_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__o21bai_1
XANTENNA__06820__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold359 final_design.cpu.reg_window\[64\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11100__A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout806 net807 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__buf_4
XFILLER_0_1_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout817 _02095_ vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_2
X_09861_ net480 _04397_ net493 vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__o21a_1
Xfanout828 net829 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09208__C net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout839 net840 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_4
X_08812_ _03759_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__nand2_1
Xhold1004 final_design.cpu.reg_window\[424\] vssd1 vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
X_09792_ net544 net543 net541 net540 net454 net463 vssd1 vssd1 vccd1 vccd1 _04711_
+ sky130_fd_sc_hd__mux4_1
Xhold1015 final_design.cpu.reg_window\[275\] vssd1 vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 final_design.cpu.reg_window\[384\] vssd1 vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07724__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__A _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08743_ _03693_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__inv_2
Xhold1037 final_design.cpu.reg_window\[425\] vssd1 vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 final_design.cpu.reg_window\[301\] vssd1 vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07128__A1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1059 final_design.cpu.reg_window\[105\] vssd1 vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout181_A _06074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12121__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09999__X _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08674_ _03622_ _03623_ _03624_ _03618_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__o211a_1
X_07625_ _02573_ _02575_ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_159_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11880__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1090_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout446_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07556_ _01469_ _02094_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__nand2_1
XANTENNA__12424__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06507_ _01377_ net1051 net1007 net1004 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__or4_2
XFILLER_0_9_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11632__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10435__B2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07487_ _02215_ _02437_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout613_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09226_ _03521_ _03640_ _03520_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_146_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09053__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09157_ net551 net549 net548 net547 net458 net467 vssd1 vssd1 vccd1 vccd1 _04076_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09425__A_N _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08108_ final_design.cpu.reg_window\[716\] final_design.cpu.reg_window\[748\] net847
+ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__mux2_1
XANTENNA__09239__X _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08290__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09088_ _02300_ _02433_ net628 vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08039_ net725 _02989_ net888 vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08239__S0 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold860 final_design.cpu.reg_window\[359\] vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 final_design.cpu.reg_window\[601\] vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 final_design.cpu.reg_window\[215\] vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ _01387_ _05772_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__and2_1
Xhold893 final_design.cpu.reg_window\[304\] vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ net83 _04191_ net84 vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07634__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07206__Y _02157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11952_ _06153_ net291 net410 net2174 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__a22o_1
XANTENNA__09134__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10903_ net82 _05610_ _05632_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_28_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11871__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11883_ net679 _06116_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__nand2_2
XFILLER_0_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13622_ clknet_leaf_124_clk _00853_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[610\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10834_ net78 net1055 vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06774__A _01718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12415__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10426__B2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13553_ clknet_leaf_105_clk _00784_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[541\]
+ sky130_fd_sc_hd__dfrtp_1
X_10765_ _05438_ _05457_ _05478_ _05498_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__nand4_1
XFILLER_0_67_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09292__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12504_ _06166_ net344 net327 net1875 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13484_ clknet_leaf_118_clk _00715_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[472\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10696_ net39 _05435_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12435_ net2050 net227 net337 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07809__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09296__S _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13004__RESET_B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12366_ net1683 net242 net272 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__mux2_1
XANTENNA__06713__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14105_ clknet_leaf_82_clk _01302_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11317_ net2547 net317 _06011_ net434 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12297_ net1689 net232 net367 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__mux2_1
X_14036_ clknet_leaf_51_clk _00006_ net1155 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11248_ net598 _05949_ _05950_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__and3_1
XANTENNA__12351__B2 final_design.cpu.reg_window\[820\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12450__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ _04846_ _05143_ net600 _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__o211a_2
XANTENNA__09325__A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11574__B net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12103__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10665__A1 _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11862__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07410_ net752 net675 net703 _01496_ _02360_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__o221a_2
XANTENNA__11590__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08390_ final_design.cpu.reg_window\[838\] final_design.cpu.reg_window\[870\] net830
+ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__mux2_1
XANTENNA__12406__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11614__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07341_ _02288_ _02289_ _02290_ _02291_ net783 net793 vssd1 vssd1 vccd1 vccd1 _02292_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_169_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06716__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10968__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07272_ final_design.cpu.reg_window\[134\] final_design.cpu.reg_window\[166\] net914
+ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09011_ _03735_ _03741_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold101 net103 vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 final_design.cpu.reg_window\[218\] vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 final_design.VGA_data_control.data_to_VGA\[17\] vssd1 vssd1 vccd1 vccd1 net1476
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 final_design.VGA_data_control.ready_data\[16\] vssd1 vssd1 vccd1 vccd1 net1487
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12590__B2 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold145 final_design.cpu.reg_window\[199\] vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold156 final_design.VGA_data_control.ready_data\[27\] vssd1 vssd1 vccd1 vccd1 net1509
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 final_design.cpu.reg_window\[722\] vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 final_design.VGA_data_control.ready_data\[25\] vssd1 vssd1 vccd1 vccd1 net1531
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _03423_ _04087_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__nand2_1
Xhold189 final_design.VGA_data_control.ready_data\[5\] vssd1 vssd1 vccd1 vccd1 net1542
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _03627_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__buf_4
XFILLER_0_111_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout614 net615 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout396_A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__buf_2
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 _06192_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__buf_4
Xfanout647 net648 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__buf_4
X_09844_ _04761_ _04762_ _04760_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__a21oi_1
Xfanout658 _05849_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_2
XANTENNA__10353__B1 _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1103_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 _02511_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_4
X_09775_ net497 _04693_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout563_A _06238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06987_ net900 _01930_ _01936_ _01923_ _01924_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a32o_4
XFILLER_0_38_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout184_X net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ final_design.CPU_instr_adr\[17\] _01909_ vssd1 vssd1 vccd1 vccd1 _03677_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08657_ net613 _02635_ _02611_ _01453_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__o211a_1
XANTENNA__11853__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09889__B net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout730_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout828_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06955__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07608_ final_design.cpu.reg_window\[605\] final_design.cpu.reg_window\[637\] net880
+ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__mux2_1
XANTENNA__08285__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08588_ final_design.cpu.reg_window\[960\] final_design.cpu.reg_window\[992\] net862
+ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07539_ final_design.cpu.reg_window\[863\] final_design.cpu.reg_window\[895\] net926
+ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09813__A3 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10550_ final_design.CPU_instr_adr\[5\] _05277_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_4_10__f_clk_X clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09209_ _02868_ _02900_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10481_ _05221_ _05228_ _05230_ _05172_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a31o_1
XANTENNA__10844__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12220_ net571 _06148_ net507 net376 net1885 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__a32o_1
XFILLER_0_122_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11659__B net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07588__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ _06017_ net2534 net387 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__mux2_1
XANTENNA__09982__C1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11102_ final_design.CPU_instr_adr\[31\] _05822_ net1067 vssd1 vssd1 vccd1 vccd1
+ _05823_ sky130_fd_sc_hd__mux2_1
X_12082_ net2464 net394 net503 _06011_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__a22o_1
Xhold690 final_design.cpu.reg_window\[329\] vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11675__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ _05673_ _05753_ _05754_ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a31oi_4
XANTENNA__09734__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07364__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ net1326 _00215_ net1224 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11935_ _06136_ net281 net410 net2024 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__a22o_1
X_14240__1305 vssd1 vssd1 vccd1 vccd1 _14240__1305/HI net1305 sky130_fd_sc_hd__conb_1
XFILLER_0_157_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11866_ net2450 net520 _06243_ net427 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__a22o_1
X_13605_ clknet_leaf_4_clk _00836_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[593\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10817_ _05530_ _05533_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11797_ net2568 net414 _06235_ net436 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_60_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13536_ clknet_leaf_37_clk _00767_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[524\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07276__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ net74 net1056 vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__and2_1
XANTENNA__07815__A2 _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13467_ clknet_leaf_154_clk _00698_ net1117 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[455\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12445__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10679_ _05419_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11202__X _05910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07539__S net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12418_ final_design.cpu.reg_window\[885\] net342 vssd1 vssd1 vccd1 vccd1 _06280_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12021__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13398_ clknet_leaf_128_clk _00629_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[386\]
+ sky130_fd_sc_hd__dfrtp_1
X_12349_ net2311 net360 net343 _05997_ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10583__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11127__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06910_ _01857_ _01858_ _01859_ _01860_ net774 net795 vssd1 vssd1 vccd1 vccd1 _01861_
+ sky130_fd_sc_hd__mux4_1
X_14019_ clknet_leaf_6_clk _01250_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1007\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14044__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07890_ final_design.cpu.reg_window\[279\] final_design.cpu.reg_window\[311\] net852
+ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06841_ final_design.cpu.reg_window\[276\] final_design.cpu.reg_window\[308\] net953
+ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10886__B2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09560_ _04356_ _04358_ _04390_ _04424_ _04478_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__o2111a_1
XANTENNA__12088__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06772_ _01718_ _01722_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08511_ _03458_ _03459_ _03460_ _03461_ net693 net712 vssd1 vssd1 vccd1 vccd1 _03462_
+ sky130_fd_sc_hd__mux4_1
X_09491_ _04408_ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_19_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08442_ final_design.cpu.reg_window\[260\] final_design.cpu.reg_window\[292\] net859
+ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10648__B final_design.VGA_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08373_ net607 _03321_ _03297_ _02211_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_173_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07324_ _02271_ _02272_ _02273_ _02274_ net783 net802 vssd1 vssd1 vccd1 vccd1 _02275_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12260__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09008__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07255_ final_design.cpu.reg_window\[647\] final_design.cpu.reg_window\[679\] net937
+ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout311_A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout409_A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12012__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07186_ final_design.cpu.reg_window\[137\] final_design.cpu.reg_window\[169\] net924
+ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1220_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07665__S1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout400 net403 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_8
Xfanout411 _06252_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_4
XANTENNA_fanout778_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 net424 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07692__B _02513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout433 net436 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06589__A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11926__C net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout444 net445 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_4
Xfanout455 net456 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_4
Xfanout466 net467 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_2
X_09827_ net99 _04181_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__nand2_1
Xfanout477 net479 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_2
Xfanout488 net489 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_2
XANTENNA_fanout945_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout499 _03418_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12079__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ net451 _04675_ _04672_ net735 vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__a211o_2
X_08709_ _01359_ _01599_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__nor2_1
XANTENNA__11826__A0 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ net485 _04607_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11434__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ net435 net586 _06218_ net297 net1789 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__a32o_1
XFILLER_0_90_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout900_X net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11651_ net192 net638 vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10602_ net1474 net1046 net1016 _05346_ vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__a22o_1
XANTENNA__11054__B2 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12251__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11582_ net194 net642 vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13321_ clknet_leaf_89_clk _00552_ net1233 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[309\]
+ sky130_fd_sc_hd__dfrtp_1
X_10533_ net814 _05276_ _05280_ net975 vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__o22a_1
XFILLER_0_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_9__f_clk_X clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12003__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13252_ clknet_leaf_93_clk _00483_ net1227 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[240\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input74_A memory_size[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ _04940_ net252 vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__nor2_1
XANTENNA__11389__B net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07105__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ net573 _06131_ net509 net376 net2041 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__a32o_1
XANTENNA__11357__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13183_ clknet_leaf_134_clk _00414_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[171\]
+ sky130_fd_sc_hd__dfrtp_1
X_10395_ net813 net1016 _05179_ net1045 net2310 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__a32o_1
X_12134_ net239 net2499 net386 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09970__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11109__A2 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12306__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09707__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ net2385 net394 net502 _05884_ vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_53_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09183__B1 _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11016_ _05720_ _05722_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__nor2_1
XANTENNA__09722__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11817__A0 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ clknet_leaf_43_clk _00205_ net1150 vssd1 vssd1 vccd1 vccd1 final_design.uart.bits_received\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09486__A1 _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10749__A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12085__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11293__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ final_design.cpu.reg_window\[414\] _05845_ vssd1 vssd1 vccd1 vccd1 _06251_
+ sky130_fd_sc_hd__or2_1
XANTENNA__12490__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12898_ clknet_leaf_55_clk _00136_ net1160 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11849_ _06099_ net288 net522 net2524 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12242__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_109_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12175__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13519_ clknet_leaf_92_clk _00750_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[507\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload10 clknet_leaf_166_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_6
Xclkload21 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__clkinv_2
X_07040_ final_design.cpu.reg_window\[718\] final_design.cpu.reg_window\[750\] net935
+ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__mux2_1
Xclkload32 clknet_leaf_159_clk vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_42_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload43 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_141_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload54 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload54/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload65 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__inv_6
XFILLER_0_140_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload76 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_77_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload87 clknet_leaf_139_clk vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_149_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload98 clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__clkinv_4
X_08991_ _03792_ _03926_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__or2_2
XFILLER_0_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07942_ net725 _02892_ net888 vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_166_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10843__A2_N net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07873_ final_design.cpu.reg_window\[724\] final_design.cpu.reg_window\[756\] net866
+ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ _04529_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__xnor2_1
X_06824_ final_design.cpu.reg_window\[917\] final_design.cpu.reg_window\[949\] net963
+ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07732__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09543_ net497 _04461_ _04231_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__a21oi_1
X_06755_ final_design.cpu.reg_window\[791\] final_design.cpu.reg_window\[823\] net919
+ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__mux2_1
XANTENNA__11808__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__A net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_A _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09477__A1 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout359_A _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ net543 net541 net540 net539 net457 net466 vssd1 vssd1 vccd1 vccd1 _04393_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06686_ _01633_ _01634_ _01635_ _01636_ net784 net802 vssd1 vssd1 vccd1 vccd1 _01637_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12481__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08425_ final_design.cpu.reg_window\[901\] final_design.cpu.reg_window\[933\] net823
+ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1170_A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout526_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08356_ _03303_ _03304_ _03305_ _03306_ net685 net706 vssd1 vssd1 vccd1 vccd1 _03307_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12233__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06872__A _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload4 clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_6
X_07307_ final_design.cpu.reg_window\[901\] final_design.cpu.reg_window\[933\] net906
+ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__mux2_1
XANTENNA__11587__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08287_ net719 _03237_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07238_ final_design.cpu.reg_window\[135\] final_design.cpu.reg_window\[167\] net916
+ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout895_A _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07169_ final_design.cpu.reg_window\[714\] final_design.cpu.reg_window\[746\] net919
+ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1223_X net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ final_design.uart.BAUD_counter\[29\] final_design.uart.BAUD_counter\[28\]
+ final_design.uart.BAUD_counter\[31\] final_design.uart.BAUD_counter\[30\] vssd1
+ vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11429__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12773__4 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__inv_2
XFILLER_0_79_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1206 net1209 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__clkbuf_2
Xfanout1217 net100 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__buf_2
Xfanout1228 net1229 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__clkbuf_4
Xfanout230 net232 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
Xfanout241 net242 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
Xfanout1239 net1256 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__buf_2
Xfanout252 net254 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07208__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout263 net265 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout285 net286 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08912__B1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 net298 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_4
X_13870_ clknet_leaf_113_clk _01101_ net1212 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[858\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07810__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07642__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12821_ net1383 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09423__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12067__A3 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12752_ final_design.VGA_adr\[5\] net808 _06383_ _06388_ _06389_ vssd1 vssd1 vccd1
+ vccd1 _01352_ sky130_fd_sc_hd__a221o_1
XANTENNA__11275__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12472__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10288__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11703_ net221 net637 vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12683_ final_design.VGA_data_control.ready_data\[29\] net1032 net987 final_design.data_from_mem\[29\]
+ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11027__A1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11634_ net429 net578 _06174_ net300 net1473 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__a32o_1
XANTENNA__12224__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11565_ net427 net573 _06138_ net303 net1560 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07877__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06454__A1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07089__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13304_ clknet_leaf_135_clk _00535_ net1167 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[292\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10516_ _05263_ _05264_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_98_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11496_ net176 net2288 net308 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13235_ clknet_leaf_32_clk _00466_ net1129 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[223\]
+ sky130_fd_sc_hd__dfrtp_1
X_10447_ net1388 net1040 _05207_ net246 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13166_ clknet_leaf_115_clk _00397_ net1204 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[154\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10378_ net21 net1036 net1019 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1
+ vccd1 _00131_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12117_ net1825 net194 net388 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13097_ clknet_leaf_89_clk _00328_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09156__A0 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12048_ net2042 net196 net399 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11582__B net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13999_ clknet_leaf_92_clk _01230_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[987\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06540_ _01464_ _01475_ _01483_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__or3_1
XFILLER_0_172_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11266__B2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13200__RESET_B net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06471_ final_design.data_from_mem\[16\] net983 _01421_ vssd1 vssd1 vccd1 vccd1 _01422_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08210_ _02000_ net616 vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__nor2_1
XANTENNA__06693__A1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11018__B2 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12215__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08383__S net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09190_ net496 _04107_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__nand2_2
XFILLER_0_90_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06692__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11569__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08141_ final_design.cpu.reg_window\[973\] final_design.cpu.reg_window\[1005\] net832
+ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload110 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 clkload110/Y sky130_fd_sc_hd__clkinvlp_4
X_08072_ _01881_ net617 vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__nor2_1
Xclkload121 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload121/Y sky130_fd_sc_hd__inv_4
XTAP_TAPCELL_ROW_116_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload132 clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 clkload132/Y sky130_fd_sc_hd__inv_6
Xclkload143 clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 clkload143/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07023_ final_design.cpu.reg_window\[398\] final_design.cpu.reg_window\[430\] net934
+ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_168_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09395__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_126_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08974_ _03676_ _03677_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1016_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold16 final_design.cpu.reg_window\[27\] vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ final_design.cpu.reg_window\[86\] final_design.cpu.reg_window\[118\] net819
+ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__mux2_1
Xhold27 final_design.cpu.reg_window\[13\] vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 final_design.reqhand.instruction\[8\] vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 _01309_ vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ final_design.cpu.reg_window\[276\] final_design.cpu.reg_window\[308\] net872
+ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
X_06807_ _01750_ _01755_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__nand2_1
XANTENNA__08370__B2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11492__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07787_ _02737_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout643_A _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09526_ _04342_ _04439_ _04441_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__o22a_1
X_06738_ net751 net893 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09457_ _04304_ _04307_ net476 vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06669_ final_design.cpu.reg_window\[602\] final_design.cpu.reg_window\[634\] net952
+ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1173_X net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout908_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12994__RESET_B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07698__A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ _03324_ _03325_ _03355_ _03357_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__o22a_1
XANTENNA__11009__B2 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12206__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ net534 net533 _02325_ net532 net460 net470 vssd1 vssd1 vccd1 vccd1 _04307_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07308__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08339_ net619 _03287_ _03288_ net538 vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_145_970 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07859__S1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12221__A3 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ net668 _03847_ net740 vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _01384_ _05154_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout898_X net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11980__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11281_ _05844_ _05978_ _05979_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__and3_1
XANTENNA__10852__A _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13020_ clknet_leaf_149_clk _00251_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10232_ _05108_ net811 _05107_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__and3b_1
XANTENNA__11667__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__B1 _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10163_ final_design.VGA_data_control.VGA_request_address\[0\] _05054_ final_design.VGA_data_control.VGA_request_address\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__a21o_1
Xfanout1003 _01414_ vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__buf_2
XFILLER_0_100_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1014 _05239_ vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09138__A0 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08041__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1025 _05166_ vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1036 net1037 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input37_A mem_adr_start[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 net1048 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__buf_4
X_10094_ final_design.VGA_data_control.h_count\[8\] final_design.VGA_data_control.h_count\[9\]
+ _05008_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__or3_1
Xfanout1058 net1060 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12288__A3 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1069 final_design.reqhand.current_client\[2\] vssd1 vssd1 vccd1 vccd1 net1069
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11683__A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13922_ clknet_leaf_14_clk _01153_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[910\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13853_ clknet_leaf_13_clk _01084_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[841\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12804_ net1386 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__clkbuf_1
X_10996_ _05721_ _05717_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__and2b_1
X_13784_ clknet_leaf_129_clk _01015_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[772\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _06374_ _06375_ _06370_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08664__A2 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06675__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12666_ _06320_ net1438 net991 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11617_ net238 net639 vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ net1453 net1012 net998 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1
+ vccd1 _01290_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10759__B1 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12212__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11420__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11548_ net223 net642 vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold508 final_design.cpu.reg_window\[900\] vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11971__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11858__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold519 final_design.cpu.reg_window\[851\] vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
X_11479_ net197 net2479 net309 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13218_ clknet_leaf_29_clk _00449_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[206\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07547__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09328__A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14198_ net1267 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XANTENNA__11184__A0 final_design.reqhand.data_from_UART\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ clknet_leaf_10_clk _00380_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[137\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 final_design.uart.BAUD_counter\[18\] vssd1 vssd1 vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 final_design.data_from_mem\[28\] vssd1 vssd1 vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12279__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07710_ net729 _02660_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__nor2_1
X_08690_ _02419_ net456 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nand2_1
XANTENNA__08378__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ final_design.cpu.reg_window\[988\] final_design.cpu.reg_window\[1020\] net875
+ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11239__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07572_ final_design.cpu.reg_window\[31\] final_design.cpu.reg_window\[63\] net841
+ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__mux2_1
X_09311_ _04222_ _04229_ _04218_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__a21o_1
X_06523_ _01466_ _01467_ _01471_ net980 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__or4_4
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09852__A1 _04153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11532__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09242_ _02994_ _03026_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__nor2_1
X_06454_ net1072 net1052 final_design.reqhand.current_client\[1\] vssd1 vssd1 vccd1
+ vccd1 _01407_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06626__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09173_ _03635_ net666 vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__or2_2
XFILLER_0_161_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12203__A3 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout224_A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08124_ final_design.cpu.reg_window\[333\] final_design.cpu.reg_window\[365\] net834
+ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__mux2_1
XANTENNA__11411__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11962__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ final_design.cpu.reg_window\[210\] final_design.cpu.reg_window\[242\] net818
+ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1133_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09368__B1 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07006_ final_design.cpu.reg_window\[975\] final_design.cpu.reg_window\[1007\] net909
+ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08266__S1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09383__A3 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ _03751_ _03895_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout760_A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_X net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ final_design.cpu.reg_window\[599\] final_design.cpu.reg_window\[631\] net828
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__mux2_1
XANTENNA__08879__C1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08888_ net632 _03832_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__nor2_1
XANTENNA__08288__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07839_ _02786_ _02787_ _02788_ _02789_ net697 net716 vssd1 vssd1 vccd1 vccd1 _02790_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _05559_ _05564_ _05581_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12427__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07920__S net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09509_ _02936_ _04426_ _04160_ _03029_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__o211ai_1
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10781_ final_design.CPU_instr_adr\[16\] _03928_ net1070 vssd1 vssd1 vccd1 vccd1
+ _05517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12520_ _06182_ net343 net327 net2519 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11650__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10453__A2 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07854__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12451_ net2035 net200 net335 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11402_ _01501_ net650 _06085_ net653 vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11402__B2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12382_ net1703 net202 net270 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09071__A2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14121_ clknet_leaf_76_clk final_design.vga.v_next_count\[1\] net1252 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_10_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11333_ net2455 net315 _06025_ net425 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__a22o_1
XANTENNA__11953__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10059__A2_N _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14052_ clknet_leaf_47_clk _00013_ net1148 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11264_ _04613_ net659 net598 _05964_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__o211a_1
XANTENNA__11397__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11166__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ net1345 _00234_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_10215_ final_design.uart.BAUD_counter\[5\] final_design.uart.BAUD_counter\[4\] _05094_
+ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__and3_1
X_11195_ _04723_ net659 net599 _05903_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__o211a_4
X_10146_ final_design.VGA_data_control.h_count\[0\] _05046_ vssd1 vssd1 vccd1 vccd1
+ final_design.vga.h_next_count\[0\] sky130_fd_sc_hd__and2b_1
X_10077_ wb_manage.curr_state\[2\] wb_manage.curr_state\[1\] vssd1 vssd1 vccd1 vccd1
+ _04994_ sky130_fd_sc_hd__nor2_2
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12130__A2 _06268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13905_ clknet_leaf_110_clk _01136_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[893\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload2_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13836_ clknet_leaf_121_clk _01067_ net1197 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[824\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07830__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09611__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10979_ net971 _05703_ _05705_ net969 vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_139_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13767_ clknet_leaf_9_clk _00998_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[755\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12448__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08637__A2 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06648__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12718_ _06355_ _06356_ _06358_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__a21o_2
XANTENNA__09330__B _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13698_ clknet_leaf_28_clk _00929_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[686\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12649_ final_design.VGA_data_control.ready_data\[12\] net1035 net990 final_design.data_from_mem\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11588__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11944__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12183__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold305 final_design.cpu.reg_window\[59\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold316 net128 vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10492__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold327 final_design.cpu.reg_window\[692\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 final_design.cpu.reg_window\[76\] vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold349 final_design.cpu.reg_window\[191\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06820__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11157__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout807 _01418_ vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_8
X_09860_ _04641_ _04778_ net471 vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout818 net820 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_4
Xfanout829 net840 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__buf_2
X_08811_ _03760_ _03761_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__and2_1
XANTENNA__09770__B1 _04687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09791_ net539 net538 net537 net536 net453 net463 vssd1 vssd1 vccd1 vccd1 _04710_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10380__B2 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1005 final_design.cpu.reg_window\[823\] vssd1 vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 final_design.cpu.reg_window\[943\] vssd1 vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11527__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08742_ net673 _01537_ final_design.CPU_instr_adr\[9\] vssd1 vssd1 vccd1 vccd1 _03693_
+ sky130_fd_sc_hd__a21oi_1
Xhold1027 final_design.cpu.reg_window\[354\] vssd1 vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12657__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1038 final_design.cpu.reg_window\[997\] vssd1 vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 final_design.cpu.reg_window\[827\] vssd1 vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08673_ _01999_ _02062_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07624_ net613 _02570_ _02546_ net561 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__o211a_1
XANTENNA__12409__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07555_ _01469_ _02094_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__and2_2
XFILLER_0_119_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11770__B net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout341_A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10667__A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06506_ final_design.data_from_mem\[4\] _01393_ net1006 net1003 vssd1 vssd1 vccd1
+ vccd1 _01457_ sky130_fd_sc_hd__and4_1
XFILLER_0_146_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11632__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10435__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07486_ _02242_ _02436_ _02241_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10386__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09225_ _03262_ _03293_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__and2_1
X_06437_ net35 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout606_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout227_X net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09156_ net555 net554 net553 net552 net458 net467 vssd1 vssd1 vccd1 vccd1 _04075_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06880__A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08107_ _03054_ _03055_ _03056_ _03057_ net687 net708 vssd1 vssd1 vccd1 vccd1 _03058_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11935__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09087_ final_design.CPU_instr_adr\[5\] _04011_ net1050 vssd1 vssd1 vccd1 vccd1 _00216_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__08261__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_142_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07187__S net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08038_ _02985_ _02986_ _02987_ _02988_ net683 net699 vssd1 vssd1 vccd1 vccd1 _02989_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold850 final_design.cpu.reg_window\[922\] vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout975_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08239__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold861 final_design.cpu.reg_window\[771\] vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13374__RESET_B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold872 final_design.cpu.reg_window\[879\] vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 final_design.cpu.reg_window\[249\] vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 final_design.cpu.reg_window\[316\] vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ _04918_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__inv_2
XANTENNA__12360__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ _04370_ _04773_ _04409_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10371__B2 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _06152_ net292 net411 net2148 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__a22o_1
XANTENNA__14110__Q final_design.reqhand.data_from_UART\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10902_ _05630_ _05631_ _05610_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_28_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11871__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11882_ net177 net648 net285 net521 net1907 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__a32o_1
XFILLER_0_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10833_ _04571_ net251 _04990_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__o21ai_1
X_13621_ clknet_leaf_53_clk _00852_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[609\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06774__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10426__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09150__B _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10764_ net1015 _05499_ _05500_ net1041 net1449 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__a32o_1
X_13552_ clknet_leaf_104_clk _00783_ net1204 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[540\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08047__A _01881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09292__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12503_ _06165_ net344 net327 net1938 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13483_ clknet_leaf_20_clk _00714_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[471\]
+ sky130_fd_sc_hd__dfrtp_1
X_10695_ net676 _05424_ _05434_ net977 _05433_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__o221a_1
XFILLER_0_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11900__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12434_ net1673 net241 net337 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08481__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12365_ net1778 net228 net271 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_101_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07097__S net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06802__A1 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14104_ clknet_leaf_96_clk _01301_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11316_ net656 net587 net197 vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and3_1
X_12296_ _05867_ _06260_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14035_ clknet_leaf_35_clk _01266_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1023\]
+ sky130_fd_sc_hd__dfrtp_1
X_11247_ _04639_ _04653_ net659 vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12351__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07825__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ net665 _05886_ _05888_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__or3_1
XANTENNA__10362__B2 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ final_design.vga.v_current_state\[0\] _05034_ _04999_ vssd1 vssd1 vccd1 vccd1
+ _05035_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_168_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_168_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10665__A2 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11590__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13819_ clknet_leaf_155_clk _01050_ net1115 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[807\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12178__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07340_ final_design.cpu.reg_window\[516\] final_design.cpu.reg_window\[548\] net941
+ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11614__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06716__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07271_ final_design.cpu.reg_window\[198\] final_design.cpu.reg_window\[230\] net914
+ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09010_ _01364_ net1049 _03943_ vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08391__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11378__B1 _06064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold102 net161 vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold113 final_design.cpu.reg_window\[195\] vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 net148 vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 net129 vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold146 final_design.VGA_data_control.ready_data\[6\] vssd1 vssd1 vccd1 vccd1 net1499
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09418__S0 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold157 net154 vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 net153 vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 final_design.cpu.reg_window\[158\] vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09912_ _04149_ _04830_ net450 vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10950__A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout604 net605 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_2
Xfanout615 _02514_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__clkbuf_4
Xfanout626 _02513_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12342__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout637 _06192_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__buf_2
X_09843_ _03230_ _04495_ net322 vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08420__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout648 _06093_ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10353__B2 final_design.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 net660 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_4
XANTENNA_fanout291_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_A _06265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09774_ net491 _04690_ _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__o21a_1
X_06986_ net900 _01930_ _01936_ _01923_ _01924_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a32oi_4
X_08725_ final_design.CPU_instr_adr\[17\] _01909_ vssd1 vssd1 vccd1 vccd1 _03676_
+ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_159_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_159_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout556_A net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_X net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ net561 _02572_ _03606_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06955__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ net723 _02551_ net732 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_1_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ final_design.cpu.reg_window\[768\] final_design.cpu.reg_window\[800\] net870
+ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout723_A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07538_ net761 _02482_ net755 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07469_ _01489_ _01495_ _01820_ _01817_ _01816_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09208_ _04126_ _04123_ net264 vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__and3b_1
X_10480_ _05228_ _05230_ _05221_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12772__3_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__B1 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09139_ net541 net540 net539 net538 net458 net466 vssd1 vssd1 vccd1 vccd1 _04058_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12150_ net197 net2433 net386 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout880_X net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ _05820_ _05821_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout978_X net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11956__A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ net2441 net392 net500 _06004_ vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__a22o_1
Xhold680 final_design.cpu.reg_window\[1010\] vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_127_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06891__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold691 final_design.cpu.reg_window\[529\] vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07645__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ _05748_ _05755_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__nand2_1
XANTENNA__12333__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09734__B1 _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11675__B net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__B2 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06643__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12097__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ net1325 _00214_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11691__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08476__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11934_ _06135_ net287 net409 net1966 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11865_ net204 net563 vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13604_ clknet_leaf_94_clk _00835_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[592\]
+ sky130_fd_sc_hd__dfrtp_1
X_10816_ net77 _05529_ _05549_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_83_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11796_ net656 net565 net197 vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_60_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07276__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13535_ clknet_leaf_133_clk _00766_ net1166 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[523\]
+ sky130_fd_sc_hd__dfrtp_1
X_10747_ _05467_ _05470_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10678_ _05406_ _05414_ _05417_ net38 vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__a31oi_2
XANTENNA__06724__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13466_ clknet_leaf_163_clk _00697_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[454\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09100__S net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12417_ _06109_ net355 net341 net2132 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__a22o_1
X_13397_ clknet_leaf_27_clk _00628_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[385\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09973__B1 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12348_ net2366 net360 net343 _05990_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12279_ net569 _06209_ net506 net368 net2165 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__a32o_1
XANTENNA__12461__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09725__A0 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ clknet_leaf_29_clk _01249_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1006\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10335__B2 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06840_ final_design.cpu.reg_window\[340\] final_design.cpu.reg_window\[372\] net955
+ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06771_ net750 net727 net672 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__a21o_2
XANTENNA__12088__A1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08510_ final_design.cpu.reg_window\[386\] final_design.cpu.reg_window\[418\] net860
+ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__mux2_1
XANTENNA__08387__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11296__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09490_ _04093_ _04340_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__or2_2
XANTENNA__08386__S net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14013__RESET_B net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08441_ final_design.cpu.reg_window\[324\] final_design.cpu.reg_window\[356\] net859
+ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08372_ _02212_ net607 vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_173_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11599__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07323_ final_design.cpu.reg_window\[388\] final_design.cpu.reg_window\[420\] net940
+ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__mux2_1
XANTENNA__11063__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12260__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07254_ final_design.cpu.reg_window\[711\] final_design.cpu.reg_window\[743\] net915
+ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
XANTENNA__06634__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07185_ final_design.cpu.reg_window\[201\] final_design.cpu.reg_window\[233\] net924
+ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout304_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1046_A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08767__A1 final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__C1 _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11771__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12371__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout401 net403 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_4
XANTENNA__12948__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout412 net415 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_8
Xfanout423 net424 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_4
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout673_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10326__B2 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 _04090_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_2
Xfanout456 _03552_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_2
X_09826_ net735 _04744_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__nor2_1
Xfanout467 _03518_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06625__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout478 net479 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_2
Xfanout489 _03454_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_2
XANTENNA__12079__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ net451 _04675_ _04672_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__a21o_1
X_06969_ final_design.cpu.reg_window\[208\] final_design.cpu.reg_window\[240\] net958
+ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout938_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ final_design.CPU_instr_adr\[28\] _01570_ vssd1 vssd1 vccd1 vccd1 _03659_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08296__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09688_ _04434_ _04606_ net471 vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09495__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _03586_ _03588_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11650_ net425 net567 _06182_ net299 net1823 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10601_ _05329_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__xor2_1
X_11581_ net438 net595 _06146_ net306 net1622 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__a32o_1
XANTENNA__09652__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10532_ net971 _05275_ _05279_ net969 vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__o22a_1
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13320_ clknet_leaf_117_clk _00551_ net1192 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[308\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13251_ clknet_leaf_6_clk _00482_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[239\]
+ sky130_fd_sc_hd__dfrtp_1
X_10463_ net2535 net1043 _05215_ net246 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__a22o_1
XANTENNA__07105__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10014__B1 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ net568 _06130_ net505 net376 net1671 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__a32o_1
XANTENNA__12554__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13182_ clknet_leaf_21_clk _00413_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[170\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input67_A mem_adr_start[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ _03613_ _04991_ _04987_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__o21ai_1
X_12133_ net226 net2525 net386 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07981__A2 _02929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12064_ net2448 net394 net502 _05876_ vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__a22o_1
XANTENNA__10317__B2 final_design.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ _05738_ _05739_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_53_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09722__A3 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout990 _06299_ vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12966_ clknet_leaf_66_clk _00204_ net1220 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09486__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ net181 net2081 net277 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11293__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12897_ clknet_leaf_87_clk _00135_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_142_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11848_ _06098_ net289 net522 net2332 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09238__A2 _04153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13477__RESET_B net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12797__28 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__inv_2
XFILLER_0_145_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12242__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12456__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11779_ net2500 net412 net281 _05911_ vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__a22o_1
XANTENNA__13406__RESET_B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13518_ clknet_leaf_114_clk _00749_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[506\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload11 clknet_leaf_167_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload22 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_6
X_13449_ clknet_leaf_89_clk _00680_ net1234 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[437\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload33 clknet_leaf_160_clk vssd1 vssd1 vccd1 vccd1 clkload33/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__09946__A0 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload44 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload44/X sky130_fd_sc_hd__clkbuf_8
Xclkload55 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 clkload55/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__12545__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload66 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload77 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__inv_8
XFILLER_0_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11753__A0 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload88 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_149_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload99 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__inv_8
XANTENNA__11596__A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12191__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ final_design.CPU_instr_adr\[15\] _03791_ final_design.CPU_instr_adr\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08241__Y _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09066__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ _02888_ _02889_ _02890_ _02891_ net682 net699 vssd1 vssd1 vccd1 vccd1 _02892_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_166_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07872_ net721 _02822_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__nor2_1
XANTENNA__06607__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ net86 _04193_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_3_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06823_ final_design.cpu.reg_window\[981\] final_design.cpu.reg_window\[1013\] net963
+ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11535__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06754_ final_design.cpu.reg_window\[855\] final_design.cpu.reg_window\[887\] net918
+ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09542_ net485 _04366_ _04460_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09513__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06629__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09477__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12928__Q net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09473_ _04171_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__nand2_1
X_06685_ final_design.cpu.reg_window\[409\] final_design.cpu.reg_window\[441\] net944
+ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout254_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_90_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08424_ final_design.cpu.reg_window\[965\] final_design.cpu.reg_window\[997\] net823
+ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08355_ final_design.cpu.reg_window\[135\] final_design.cpu.reg_window\[167\] net833
+ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_9__f_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__12366__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12233__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_A net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1163_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout519_A _06259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ final_design.cpu.reg_window\[965\] final_design.cpu.reg_window\[997\] net906
+ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload5 clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08286_ _03233_ _03234_ _03235_ _03236_ net688 net709 vssd1 vssd1 vccd1 vccd1 _03237_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11992__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07237_ final_design.cpu.reg_window\[199\] final_design.cpu.reg_window\[231\] net916
+ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_X net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12536__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09937__B1 _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07099__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07168_ net759 _02118_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout888_A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__C1 _01750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07099_ _02046_ _02047_ _02048_ _02049_ net779 net800 vssd1 vssd1 vccd1 vccd1 _02050_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07195__S net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1207 net1209 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__clkbuf_4
Xfanout220 _05921_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_2
Xfanout1218 net1256 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__buf_4
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1229 net1239 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__buf_2
Xfanout231 net232 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_2
Xfanout242 _05875_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_2
Xfanout253 net255 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07208__B _02157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout264 net265 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08373__C1 _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 net277 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_4
Xfanout286 net287 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_4
Xfanout297 net298 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_8
X_09809_ _04727_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11445__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ net1372 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09423__B _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12751_ _06351_ _06372_ net967 _05058_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__and4b_1
XFILLER_0_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_81_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11702_ net569 net420 _06209_ net295 net1963 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__a32o_1
X_12682_ _06328_ net2169 net991 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11633_ net207 net639 vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__and2_1
XANTENNA__12224__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12129__X _06268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08979__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08523__S0 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11564_ net209 net642 vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11983__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13303_ clknet_leaf_143_clk _00534_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[291\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10515_ _05250_ _05260_ _05262_ net61 vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__a31o_1
XANTENNA__07651__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11495_ net178 net2351 net308 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12527__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09928__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13234_ clknet_leaf_39_clk _00465_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[222\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10446_ _02863_ net601 vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10377_ net20 net1038 net1021 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1
+ vccd1 _00130_ sky130_fd_sc_hd__a22o_1
X_13165_ clknet_leaf_103_clk _00396_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[153\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08600__B1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ net2051 net196 net391 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13096_ clknet_leaf_125_clk _00327_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09156__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12047_ net1692 net197 net398 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12160__A0 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11863__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07405__Y _02356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13998_ clknet_leaf_114_clk _01229_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[986\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08116__C1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12949_ clknet_leaf_55_clk _00187_ net1160 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11266__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12463__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_72_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06470_ final_design.reqhand.instruction\[16\] net982 vssd1 vssd1 vccd1 vccd1 _01421_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_157_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12186__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08140_ final_design.cpu.reg_window\[781\] final_design.cpu.reg_window\[813\] net832
+ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__mux2_1
XANTENNA__07140__Y _02091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11974__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08071_ net888 _03021_ _03010_ _03009_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__o2bb2a_4
Xclkload100 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 clkload100/Y sky130_fd_sc_hd__bufinv_16
Xclkload111 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 clkload111/Y sky130_fd_sc_hd__clkinv_2
Xclkload122 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 clkload122/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_116_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12518__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07022_ final_design.cpu.reg_window\[462\] final_design.cpu.reg_window\[494\] net935
+ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__mux2_1
Xclkload133 clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 clkload133/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload144 clknet_leaf_80_clk vssd1 vssd1 vccd1 vccd1 clkload144/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__06912__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_168_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11726__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07945__A2 _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ final_design.CPU_instr_adr\[18\] net1027 _03908_ _03910_ vssd1 vssd1 vccd1
+ vccd1 _00229_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold17 final_design.cpu.reg_window\[28\] vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 net118 vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ net717 _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__nor2_1
Xhold39 final_design.cpu.reg_window\[7\] vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A _06295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07743__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07253__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09524__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ final_design.cpu.reg_window\[340\] final_design.cpu.reg_window\[372\] net873
+ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout469_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06806_ _01750_ _01755_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07786_ _02734_ _02736_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__nor2_1
XANTENNA__13399__RESET_B net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09525_ _04116_ _04443_ _04442_ net321 vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__a2bb2o_1
X_06737_ net891 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__inv_2
XANTENNA__12454__A1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10465__A0 final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_63_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout636_A _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06668_ net763 _01618_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__or2_1
XANTENNA__08574__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ net476 _04302_ _04374_ net320 vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08407_ _03355_ _03357_ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__or2_2
XFILLER_0_109_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12096__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06599_ final_design.cpu.reg_window\[476\] final_design.cpu.reg_window\[508\] net954
+ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout803_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ net490 _04305_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07308__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08338_ net605 _03287_ _03263_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__o21a_1
XANTENNA__09622__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11965__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08269_ final_design.cpu.reg_window\[586\] final_design.cpu.reg_window\[618\] net837
+ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10300_ final_design.VGA_data_control.data_to_VGA\[11\] final_design.VGA_data_control.data_to_VGA\[10\]
+ final_design.VGA_data_control.data_to_VGA\[9\] final_design.VGA_data_control.data_to_VGA\[8\]
+ net1063 net1062 vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09258__X _04177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12509__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ _04681_ _04696_ net659 vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__a21o_1
XANTENNA__06822__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10852__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ final_design.uart.BAUD_counter\[11\] final_design.uart.BAUD_counter\[10\]
+ _05104_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06819__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__A1 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10162_ final_design.VGA_data_control.VGA_request_address\[0\] _05054_ _05056_ vssd1
+ vssd1 vccd1 vccd1 final_design.vga.h_next_count\[6\] sky130_fd_sc_hd__o21a_1
XANTENNA__11018__A2_N net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07219__A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1004 _01413_ vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_2
Xfanout1015 net1017 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09138__A1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14113__Q final_design.reqhand.data_from_UART\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1026 net1027 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10093_ final_design.VGA_data_control.h_count\[8\] final_design.VGA_data_control.h_count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__nor2_1
Xfanout1037 _05169_ vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1048 _04994_ vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12142__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 net1060 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__buf_1
X_13921_ clknet_leaf_155_clk _01152_ net1113 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[909\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11683__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13852_ clknet_leaf_153_clk _01083_ net1118 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[840\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09153__B net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12803_ net1376 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13783_ clknet_leaf_137_clk _01014_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[771\]
+ sky130_fd_sc_hd__dfrtp_1
X_10995_ net86 _05698_ _05720_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__a21o_1
XANTENNA__11903__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12734_ _06364_ _06367_ _06368_ final_design.VGA_data_control.v_count\[0\] vssd1
+ vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_48_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08484__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12665_ final_design.VGA_data_control.ready_data\[20\] net1032 net987 final_design.data_from_mem\[20\]
+ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11616_ net568 net420 _06165_ net299 net1607 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_137_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12596_ net1734 net1011 net997 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1
+ vccd1 _01289_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11547_ net2543 net305 _06129_ net423 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07828__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold509 final_design.cpu.reg_window\[977\] vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06732__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11858__B net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11478_ net198 net647 vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_74_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11708__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09377__A1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13217_ clknet_leaf_158_clk _00448_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[205\]
+ sky130_fd_sc_hd__dfrtp_1
X_10429_ _03129_ _05190_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__nor2_1
X_14197_ net1266 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XANTENNA__11184__A1 final_design.data_from_mem\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ clknet_leaf_148_clk _00379_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[136\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10931__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10931__B2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ clknet_leaf_144_clk _00310_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[67\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1209 final_design.CPU_instr_adr\[30\] vssd1 vssd1 vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07640_ final_design.cpu.reg_window\[796\] final_design.cpu.reg_window\[828\] net874
+ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__mux2_1
XANTENNA__09631__X _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire225_X net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11239__A2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07571_ final_design.cpu.reg_window\[95\] final_design.cpu.reg_window\[127\] net841
+ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_45_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk
+ sky130_fd_sc_hd__clkbuf_8
X_06522_ _01466_ _01467_ _01471_ net980 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__nor4_1
XANTENNA__11813__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09310_ _04226_ _04228_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__nand2_1
XANTENNA__07799__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06453_ _01405_ _01406_ _01396_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__o21ai_1
X_09241_ _04159_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09172_ _03635_ net666 vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08123_ final_design.cpu.reg_window\[397\] final_design.cpu.reg_window\[429\] net831
+ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__mux2_1
XANTENNA__11947__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout217_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08054_ final_design.cpu.reg_window\[18\] final_design.cpu.reg_window\[50\] net818
+ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09519__A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06642__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09368__A1 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12781__12 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__inv_2
XFILLER_0_114_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07005_ final_design.cpu.reg_window\[783\] final_design.cpu.reg_window\[815\] net909
+ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07379__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1126_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11784__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _03671_ _03672_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__nand2_1
X_07907_ final_design.cpu.reg_window\[663\] final_design.cpu.reg_window\[695\] net828
+ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__mux2_1
XANTENNA__12675__B2 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ _01600_ _01601_ _02472_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13509__RESET_B net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07838_ final_design.cpu.reg_window\[917\] final_design.cpu.reg_window\[949\] net884
+ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout920_A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ final_design.cpu.reg_window\[856\] final_design.cpu.reg_window\[888\] net869
+ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09508_ _02934_ _03587_ _04426_ _03029_ _02932_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__a311o_1
XFILLER_0_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10780_ _05514_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__and2_1
XANTENNA__07303__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09439_ _04191_ _04357_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__nand2_1
XANTENNA__07854__A1 _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12450_ net1743 net202 net335 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11938__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11401_ final_design.data_from_mem\[31\] net236 net234 vssd1 vssd1 vccd1 vccd1 _06085_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11402__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12381_ net1997 net204 net270 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14120_ clknet_leaf_76_clk final_design.vga.v_next_count\[0\] net1252 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.v_count\[0\] sky130_fd_sc_hd__dfrtp_4
X_11332_ net654 net567 net194 vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__and3_1
XFILLER_0_162_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14051_ clknet_leaf_48_clk _00012_ net1148 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11263_ net651 _05960_ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_91_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11166__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ net1344 _00233_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10214_ final_design.uart.BAUD_counter\[3\] final_design.uart.BAUD_counter\[4\] _05093_
+ final_design.uart.BAUD_counter\[5\] vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11194_ net663 _05900_ _05902_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10145_ _05016_ _05045_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__or2_1
XANTENNA__08479__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07383__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13932__RESET_B net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ net813 _04988_ _04992_ _01373_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__a211oi_1
XANTENNA__09531__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13904_ clknet_leaf_112_clk _01135_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[892\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ clknet_leaf_20_clk _01066_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[823\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_67_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06727__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13766_ clknet_leaf_171_clk _00997_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[754\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10978_ final_design.CPU_instr_adr\[25\] _03854_ net1072 vssd1 vssd1 vccd1 vccd1
+ _05705_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09834__A2 _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07412__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12717_ _06347_ _06357_ _06349_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06648__A2 _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13697_ clknet_leaf_159_clk _00928_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[685\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12648_ _06311_ net1397 net993 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11929__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Left_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12579_ net1443 _06294_ _06286_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11588__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 final_design.VGA_data_control.data_to_VGA\[0\] vssd1 vssd1 vccd1 vccd1 net1659
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 final_design.cpu.reg_window\[515\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold328 final_design.cpu.reg_window\[41\] vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold339 final_design.cpu.reg_window\[532\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
X_14249_ net1314 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11157__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12354__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout808 _06333_ vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout819 net820 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_4
X_08810_ final_design.CPU_instr_adr\[21\] _01788_ vssd1 vssd1 vccd1 vccd1 _03761_
+ sky130_fd_sc_hd__or2_1
X_09790_ net492 _04607_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__nand2_1
XANTENNA__06584__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1006 final_design.cpu.reg_window\[826\] vssd1 vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_163_Left_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07146__X _02097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1017 final_design.cpu.reg_window\[352\] vssd1 vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ _03690_ _03691_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__nor2_1
Xhold1028 final_design.cpu.reg_window\[431\] vssd1 vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12657__B2 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1039 final_design.cpu.reg_window\[437\] vssd1 vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13602__RESET_B net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08672_ _01501_ _01505_ _01537_ _02028_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__or4_1
XANTENNA__11081__A_N net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07623_ _01536_ _02572_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11880__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07554_ net530 _02504_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10667__B final_design.VGA_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06505_ _01454_ _01455_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__nand2_1
X_07485_ _02269_ _02434_ _02268_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_36_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11632__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10840__A0 final_design.CPU_instr_adr\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1076_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_172_Left_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09224_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__inv_2
X_06436_ net1064 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07049__C1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12374__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ _04054_ net321 vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout501_A _06264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1243_A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__A1 _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08106_ final_design.cpu.reg_window\[908\] final_design.cpu.reg_window\[940\] net847
+ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08261__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09086_ net261 _04009_ _04010_ _04007_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_115_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08037_ final_design.cpu.reg_window\[531\] final_design.cpu.reg_window\[563\] net825
+ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1031_X net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold840 final_design.cpu.reg_window\[265\] vssd1 vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12345__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold851 final_design.cpu.reg_window\[268\] vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 final_design.cpu.reg_window\[676\] vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold873 final_design.cpu.reg_window\[403\] vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 final_design.cpu.reg_window\[108\] vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold895 final_design.cpu.reg_window\[541\] vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_X net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09988_ _02737_ _04165_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08939_ final_design.CPU_instr_adr\[22\] net1028 _03876_ _03880_ vssd1 vssd1 vccd1
+ vccd1 _00233_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ _06151_ net291 net410 net2276 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__a22o_1
XANTENNA__11320__A1 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09271__X _04190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__S net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ net82 net1060 vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__or2_1
XANTENNA__09712__A _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11871__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout923_X net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ _06115_ net286 net521 net1980 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11453__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13620_ clknet_leaf_103_clk _00851_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[608\]
+ sky130_fd_sc_hd__dfrtp_1
X_10832_ _05564_ _05565_ net110 net1041 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_45_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07232__A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13551_ clknet_leaf_93_clk _00782_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[539\]
+ sky130_fd_sc_hd__dfrtp_1
X_10763_ _05477_ _05481_ _05498_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09292__A3 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12502_ _06164_ net353 net329 net1809 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10831__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input97_A memory_size[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ clknet_leaf_2_clk _00713_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[470\]
+ sky130_fd_sc_hd__dfrtp_1
X_10694_ net1066 _05430_ net1013 final_design.CPU_instr_adr\[12\] vssd1 vssd1 vccd1
+ vccd1 _05434_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_54_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12433_ net1644 net229 net336 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__mux2_1
XANTENNA__11387__A1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12364_ net2093 net231 net272 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14103_ clknet_leaf_83_clk _01300_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11315_ _04953_ net660 net599 _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__o211a_2
XFILLER_0_50_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12295_ net580 _06225_ net511 net369 net1661 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__a32o_1
XANTENNA__08998__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14034_ clknet_leaf_39_clk _01265_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1022\]
+ sky130_fd_sc_hd__dfrtp_1
X_11246_ net651 _05943_ _05948_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11177_ final_design.data_from_mem\[4\] net252 _05855_ _05887_ vssd1 vssd1 vccd1
+ vccd1 _05888_ sky130_fd_sc_hd__o211a_1
X_10128_ final_design.vga.v_current_state\[1\] _04997_ vssd1 vssd1 vccd1 vccd1 _05034_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__08002__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12639__B2 final_design.data_from_mem\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10059_ _04571_ _04573_ _04632_ _04634_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07841__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12459__S net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11862__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13818_ clknet_leaf_161_clk _01049_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[806\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09807__A2 _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10941__A_N _05662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07142__A _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13749_ clknet_leaf_40_clk _00980_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[737\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11614__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07270_ net759 _02220_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12194__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11378__A1 _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07677__S0 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold103 net142 vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 net113 vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold125 net140 vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 final_design.reqhand.instruction\[1\] vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold147 final_design.cpu.reg_window\[176\] vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 net166 vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _03423_ _04148_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__or2_1
Xhold169 final_design.VGA_data_control.ready_data\[31\] vssd1 vssd1 vccd1 vccd1 net1522
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire557_X net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10950__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout605 net615 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__buf_2
Xfanout616 net620 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_4
Xfanout627 net629 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_4
X_09842_ _03230_ _04495_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout638 net639 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__buf_4
Xfanout649 net650 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10353__A2 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08951__C1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08071__A1_N net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07317__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ net477 _04406_ _04691_ net484 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__a211o_1
X_06985_ net773 _01935_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__or2_2
XFILLER_0_77_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout284_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08724_ _03673_ _03674_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__nand2_1
XANTENNA__11302__A1 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ _01566_ _02576_ _02604_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__or3_1
XANTENNA__12369__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout451_A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_A _01880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07606_ net729 _02556_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08586_ final_design.cpu.reg_window\[832\] final_design.cpu.reg_window\[864\] net870
+ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07537_ net769 _02487_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ _02406_ _02407_ _02418_ net898 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a22oi_4
XANTENNA__08582__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09207_ _02545_ _03608_ _04052_ _04125_ _03610_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__o311a_1
X_06419_ final_design.reqhand.instruction\[2\] vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07399_ final_design.cpu.reg_window\[706\] final_design.cpu.reg_window\[738\] net946
+ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1246_X net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__B2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07198__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09138_ net546 net545 net544 net543 net458 net467 vssd1 vssd1 vccd1 vccd1 _04057_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_115_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09069_ _02438_ net633 _03991_ net259 vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11100_ net92 _05802_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07926__S net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12080_ net566 _05997_ net505 net392 net1705 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__a32o_1
XANTENNA__06891__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 final_design.cpu.reg_window\[1023\] vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08611__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 final_design.cpu.reg_window\[148\] vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold692 final_design.cpu.reg_window\[282\] vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__A1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11031_ _05729_ _05747_ _05752_ _05732_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11675__C net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06643__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ net1324 _00213_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07661__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11691__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ _06134_ net284 net409 net2390 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07233__Y _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11864_ net2264 net523 _06242_ net437 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__a22o_1
XANTENNA__08058__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13603_ clknet_leaf_1_clk _00834_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[591\]
+ sky130_fd_sc_hd__dfrtp_1
X_10815_ _05547_ _05548_ _05529_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_138_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11795_ net2508 net412 _06234_ net426 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__a22o_1
XANTENNA__11911__S net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13534_ clknet_leaf_18_clk _00765_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[522\]
+ sky130_fd_sc_hd__dfrtp_1
X_10746_ net735 _04509_ net255 _04990_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_153_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08345__X _03296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09670__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13465_ clknet_leaf_165_clk _00696_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[453\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10677_ net38 _05406_ _05414_ _05417_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__nand4_1
XFILLER_0_129_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12557__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12416_ net200 net563 net500 net340 net1830 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__a32o_1
XANTENNA__12021__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13396_ clknet_leaf_141_clk _00627_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[384\]
+ sky130_fd_sc_hd__dfrtp_1
X_12347_ net2473 net362 net358 _05981_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10583__A2 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12278_ net582 _06208_ net513 net369 net1761 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__a32o_1
X_14017_ clknet_leaf_158_clk _01248_ net1113 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1005\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09725__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _04766_ net659 net598 _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11532__A1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06770_ final_design.data_from_mem\[23\] net981 _01719_ vssd1 vssd1 vccd1 vccd1 _01721_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__07571__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08387__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12189__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08440_ _03387_ _03389_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_19_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08371_ net607 _03321_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11599__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11821__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07322_ final_design.cpu.reg_window\[452\] final_design.cpu.reg_window\[484\] net940
+ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08464__B2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06915__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07898__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07253_ _02200_ _02201_ _02202_ _02203_ net777 net797 vssd1 vssd1 vccd1 vccd1 _02204_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12548__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07184_ _02131_ _02132_ _02133_ _02134_ net780 net799 vssd1 vssd1 vccd1 vccd1 _02135_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12012__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1039_A _05168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07746__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09716__A1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 net403 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_4
Xfanout413 net415 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_4
XFILLER_0_100_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout424 _05877_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_4
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1206_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08924__C1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 net447 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 net461 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_4
X_09825_ _04737_ _04740_ _04743_ net451 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a22o_2
Xfanout468 net470 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__buf_2
XANTENNA__06625__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 net482 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout666_A _03649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout287_X net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12988__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ _03198_ _04674_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09533__Y _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08577__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06886__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ final_design.cpu.reg_window\[16\] final_design.cpu.reg_window\[48\] net958
+ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__mux2_1
XANTENNA__09262__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ _03656_ _03657_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__and2b_1
XFILLER_0_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12099__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ net548 net547 net546 net545 net453 net462 vssd1 vssd1 vccd1 vccd1 _04606_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout833_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06899_ net894 _01831_ _01837_ _01843_ _01849_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__o32a_4
XFILLER_0_68_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08638_ _03586_ _03588_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_81_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_0__f_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ net612 _03514_ _03516_ _02390_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__o211a_2
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ _05343_ _05344_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11580_ net600 net196 net645 vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10531_ _05277_ _05278_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12539__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13250_ clknet_leaf_28_clk _00481_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[238\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12003__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10462_ _02540_ net601 vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12201_ _06129_ net502 net379 net2215 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ clknet_leaf_10_clk _00412_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[169\]
+ sky130_fd_sc_hd__dfrtp_1
X_10393_ net813 net1016 _05178_ net1047 net1413 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__a32o_1
XANTENNA__06769__A1 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07966__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09437__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ net242 net2467 net386 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09707__A1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12063_ _05865_ net581 net512 net393 net1909 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__a32o_1
XANTENNA__10317__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11514__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11014_ net86 net1059 net87 vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_53_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11906__S net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout991 _06297_ vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09172__A _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12965_ clknet_leaf_66_clk _00203_ net1220 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11916_ net182 net2114 net277 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ clknet_leaf_87_clk _00134_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_16_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12490__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09891__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11847_ _06097_ net290 net522 net2380 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11778_ net2505 net412 net281 _05905_ vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13517_ clknet_leaf_139_clk _00748_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[505\]
+ sky130_fd_sc_hd__dfrtp_1
X_10729_ _05465_ _05466_ _05446_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__o21a_1
XANTENNA__07654__C1 _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload12 clknet_leaf_168_clk vssd1 vssd1 vccd1 vccd1 clkload12/X sky130_fd_sc_hd__clkbuf_4
X_13448_ clknet_leaf_117_clk _00679_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[436\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload23 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__inv_6
XFILLER_0_141_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13446__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload34 clknet_leaf_161_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_8
XANTENNA__11202__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09946__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload45 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload56 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__bufinv_16
Xclkload67 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13379_ clknet_leaf_4_clk _00610_ net1096 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[367\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_77_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload78 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07566__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload89 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11596__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09159__C1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ final_design.cpu.reg_window\[534\] final_design.cpu.reg_window\[566\] net819
+ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_11__f_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08057__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11505__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08906__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ _02818_ _02819_ _02820_ _02821_ net695 net712 vssd1 vssd1 vccd1 vccd1 _02822_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06607__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ net733 _04513_ _04527_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__or3_4
XANTENNA__11816__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ final_design.cpu.reg_window\[789\] final_design.cpu.reg_window\[821\] net964
+ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__mux2_1
XANTENNA__12060__X _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09082__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ net483 _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06753_ net760 _01697_ net755 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__o21a_1
XANTENNA__11808__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09477__A3 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09472_ _02609_ _04167_ _04170_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__nand3_1
X_06684_ final_design.cpu.reg_window\[473\] final_design.cpu.reg_window\[505\] net944
+ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__mux2_1
XANTENNA__12481__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08423_ final_design.cpu.reg_window\[773\] final_design.cpu.reg_window\[805\] net823
+ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout247_A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06791__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08354_ final_design.cpu.reg_window\[199\] final_design.cpu.reg_window\[231\] net833
+ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07330__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07305_ final_design.cpu.reg_window\[773\] final_design.cpu.reg_window\[805\] net906
+ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload6 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload6/X sky130_fd_sc_hd__clkbuf_8
X_08285_ final_design.cpu.reg_window\[393\] final_design.cpu.reg_window\[425\] net841
+ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout414_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1156_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07236_ _02185_ _02186_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09398__C1 _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12382__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07167_ _02114_ _02115_ _02116_ _02117_ net778 net798 vssd1 vssd1 vccd1 vccd1 _02118_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07099__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07098_ final_design.cpu.reg_window\[908\] final_design.cpu.reg_window\[940\] net928
+ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout783_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07048__Y _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1111_X net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout210 _05958_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_2
Xfanout1208 net1209 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__clkbuf_2
Xfanout1219 net1224 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__buf_4
Xfanout221 _05980_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1209_X net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout232 _05858_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_2
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout950_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07176__A1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout265 _04071_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_2
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net277 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_6
X_09808_ net603 _04220_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__or2_1
Xfanout287 _06228_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_4
Xfanout298 _06194_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_4
XFILLER_0_119_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09739_ net69 net70 _04182_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__nand3_1
XFILLER_0_119_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_X clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _06351_ _06384_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__xor2_1
XANTENNA__12472__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11701_ net205 net634 vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__and2_1
XFILLER_0_166_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10288__D net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12681_ final_design.VGA_data_control.ready_data\[28\] net1032 net987 final_design.data_from_mem\[28\]
+ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__a22o_1
XANTENNA__07884__C1 _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11461__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11632_ net427 net573 _06173_ net299 net1518 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__a32o_1
XFILLER_0_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08523__S1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11563_ net428 net579 _06137_ net304 net1609 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13302_ clknet_leaf_126_clk _00533_ net1192 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[290\]
+ sky130_fd_sc_hd__dfrtp_1
X_10514_ net61 _05250_ _05260_ _05262_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__and4_1
XFILLER_0_135_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11494_ net179 net648 vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__and2_1
X_13233_ clknet_leaf_107_clk _00464_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[221\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ net1477 net1040 _05206_ net246 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13164_ clknet_leaf_123_clk _00395_ net1191 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[152\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10376_ net19 net1037 net1020 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1
+ vccd1 _00129_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12115_ net1840 net197 net390 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__mux2_1
X_13095_ clknet_leaf_7_clk _00326_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09156__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12046_ net2234 net199 net396 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09106__S net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13997_ clknet_leaf_139_clk _01228_ net1181 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[985\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12948_ clknet_leaf_55_clk _00186_ net1160 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12879_ clknet_leaf_71_clk _00117_ net1246 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07150__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08070_ _03015_ _03020_ net717 vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload101 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__inv_6
XFILLER_0_153_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload112 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 clkload112/X sky130_fd_sc_hd__clkbuf_4
Xclkload123 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload123/Y sky130_fd_sc_hd__inv_6
XFILLER_0_125_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07021_ final_design.cpu.reg_window\[270\] final_design.cpu.reg_window\[302\] net934
+ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__mux2_1
Xclkload134 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 clkload134/Y sky130_fd_sc_hd__inv_6
Xclkload145 clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 clkload145/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_140_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11726__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06602__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08972_ net256 _03909_ net1027 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06988__X _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10016__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09805__A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ _02870_ _02871_ _02872_ _02873_ net682 net704 vssd1 vssd1 vccd1 vccd1 _02874_
+ sky130_fd_sc_hd__mux4_1
Xhold18 final_design.cpu.reg_window\[20\] vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 net122 vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout197_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07854_ _01504_ _01822_ net618 vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07253__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08450__S0 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06805_ _01499_ net672 _01754_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__or3b_1
X_07785_ net610 net529 _02707_ net556 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout364_A net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__C1 _02503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09524_ net475 _04107_ _04240_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__and3_1
X_06736_ final_design.reqhand.instruction\[24\] final_design.data_from_mem\[24\] net984
+ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__mux2_4
XFILLER_0_149_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10465__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11662__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ net471 _04299_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__or2_1
XANTENNA__12377__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06667_ _01614_ _01615_ _01616_ _01617_ net786 net804 vssd1 vssd1 vccd1 vccd1 _01618_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07979__B _02929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__X _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06764__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ net610 _03352_ _03328_ _02239_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09386_ _04303_ _04304_ net476 vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07881__A2 _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06598_ final_design.cpu.reg_window\[284\] final_design.cpu.reg_window\[316\] net955
+ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08337_ _02186_ net619 vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1159_X net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07094__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08268_ final_design.cpu.reg_window\[650\] final_design.cpu.reg_window\[682\] net837
+ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout998_A _06296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ net768 _02169_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08199_ final_design.cpu.reg_window\[974\] final_design.cpu.reg_window\[1006\] net844
+ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__mux2_1
X_10230_ final_design.uart.BAUD_counter\[9\] final_design.uart.BAUD_counter\[10\]
+ _05103_ final_design.uart.BAUD_counter\[11\] vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__a31o_1
XANTENNA__08043__C1 _01850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06819__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__A2 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ final_design.VGA_data_control.VGA_request_address\[0\] _05054_ _05041_ vssd1
+ vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_7_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1005 _01413_ vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__buf_1
XANTENNA__07934__S net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1016 net1017 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_58_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09138__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1027 net1028 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10092_ final_design.VGA_data_control.VGA_request_address\[1\] final_design.VGA_data_control.VGA_request_address\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__or2_1
Xfanout1038 _05168_ vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout953_X net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1049 _01410_ vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__buf_4
X_13920_ clknet_leaf_44_clk _01151_ net1149 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[908\]
+ sky130_fd_sc_hd__dfrtp_1
X_13851_ clknet_leaf_135_clk _01082_ net1168 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[839\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12802_ net1355 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__clkbuf_1
X_13782_ clknet_leaf_126_clk _01013_ net1192 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[770\]
+ sky130_fd_sc_hd__dfrtp_1
X_10994_ _05718_ _05719_ _05698_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09846__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12733_ _06364_ _06367_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10017__D_N _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12664_ _06319_ net1423 net993 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11615_ net224 net638 vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__and2_1
XFILLER_0_143_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12595_ net2026 net1011 net997 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1
+ vccd1 _01288_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input82_X net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09449__X _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11546_ net584 net239 net644 vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__and3_1
XANTENNA__07624__A2 _02570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09168__Y _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11477_ net199 net2427 net307 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13216_ clknet_leaf_36_clk _00447_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[204\]
+ sky130_fd_sc_hd__dfrtp_1
X_10428_ net1441 net1043 _05197_ net246 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__a22o_1
X_14196_ net1265 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12381__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13147_ clknet_leaf_156_clk _00378_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[135\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ net32 net1038 net1021 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1
+ _00112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ clknet_leaf_130_clk _00309_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11219__X _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ net2417 net241 net398 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__mux2_1
XANTENNA__10695__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10695__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ net720 _02520_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__nor2_1
XANTENNA__09837__B1 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06521_ final_design.data_from_mem\[0\] final_design.data_from_mem\[1\] net1051 net1007
+ net1004 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__a2111oi_1
XPHY_EDGE_ROW_85_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11644__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10447__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12197__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06746__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09240_ _02934_ _03587_ _02932_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__a21oi_1
X_06452_ net1068 net1073 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09171_ _03628_ _03650_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08122_ final_design.cpu.reg_window\[461\] final_design.cpu.reg_window\[493\] net831
+ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06923__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08704__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08053_ final_design.cpu.reg_window\[82\] final_design.cpu.reg_window\[114\] net818
+ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07004_ final_design.cpu.reg_window\[847\] final_design.cpu.reg_window\[879\] net910
+ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12660__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1021_A _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1119_A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ final_design.CPU_instr_adr\[20\] net1027 _03891_ _03894_ vssd1 vssd1 vccd1
+ vccd1 _00231_ sky130_fd_sc_hd__a22o_1
XANTENNA__11784__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12124__A1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ final_design.cpu.reg_window\[727\] final_design.cpu.reg_window\[759\] net828
+ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08879__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ _01600_ _01601_ _02472_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__nand3_1
XFILLER_0_99_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07837_ final_design.cpu.reg_window\[981\] final_design.cpu.reg_window\[1013\] net885
+ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__mux2_1
XANTENNA__07551__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07768_ net721 _02712_ net731 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__o21a_1
XANTENNA__12427__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09507_ _03590_ _04143_ _04157_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06719_ final_design.cpu.reg_window\[280\] final_design.cpu.reg_window\[312\] net949
+ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07303__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout913_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ final_design.cpu.reg_window\[91\] final_design.cpu.reg_window\[123\] net881
+ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09438_ net82 _04190_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09369_ _04194_ _04287_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11400_ net746 _03803_ _06083_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12380_ net1970 net221 net273 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__mux2_1
XANTENNA__09461__D1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08614__A net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11331_ net663 _06022_ _06023_ net598 vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__o211a_4
XFILLER_0_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ clknet_leaf_48_clk _00011_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11262_ _02000_ net649 _05962_ net661 vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_132_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13001_ net1343 _00232_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_10213_ net2551 _05094_ _05096_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__a21oi_1
X_11193_ final_design.data_from_mem\[6\] net254 _05855_ _05901_ vssd1 vssd1 vccd1
+ vccd1 _05902_ sky130_fd_sc_hd__o211a_1
XANTENNA__10374__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07664__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A mem_adr_start[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _01389_ _05044_ _05042_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10075_ net2559 _01372_ wb_manage.curr_state\[0\] _04992_ vssd1 vssd1 vccd1 vccd1
+ _00005_ sky130_fd_sc_hd__a22o_1
XANTENNA__08414__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09732__X _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13903_ clknet_leaf_90_clk _01134_ net1233 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[891\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11874__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13972__RESET_B net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13834_ clknet_leaf_164_clk _01065_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[822\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08495__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13765_ clknet_leaf_164_clk _00996_ net1085 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[753\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11626__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ final_design.CPU_instr_adr\[25\] _05703_ net1067 vssd1 vssd1 vccd1 vccd1
+ _05704_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06728__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11215__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12716_ final_design.VGA_data_control.v_count\[3\] _06348_ _06350_ vssd1 vssd1 vccd1
+ vccd1 _06357_ sky130_fd_sc_hd__o21ai_1
X_13696_ clknet_leaf_44_clk _00927_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[684\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12647_ final_design.VGA_data_control.ready_data\[11\] net1034 net989 final_design.data_from_mem\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12578_ net1065 net35 vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10773__B _04697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11529_ net1599 net189 net526 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold307 final_design.cpu.reg_window\[462\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold318 final_design.cpu.reg_window\[677\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ net1313 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
Xhold329 final_design.reqhand.instruction\[3\] vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09907__X _04826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14179_ clknet_leaf_73_clk _01353_ net1246 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08530__Y _03481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14007__RESET_B net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06979__A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout809 net810 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07574__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09770__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ final_design.CPU_instr_adr\[10\] _02128_ vssd1 vssd1 vccd1 vccd1 _03691_
+ sky130_fd_sc_hd__nor2_1
Xhold1007 final_design.cpu.reg_window\[679\] vssd1 vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 final_design.cpu.reg_window\[364\] vssd1 vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12657__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1029 final_design.cpu.reg_window\[480\] vssd1 vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10668__A1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08671_ _01568_ _01598_ _01628_ _01659_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__or4_1
XFILLER_0_139_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11824__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07622_ net626 _02570_ _02571_ net561 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12409__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07553_ net749 _01497_ _01502_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_75_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06504_ net1053 net1006 net1003 _01374_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a31o_1
XFILLER_0_159_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07484_ _02270_ _02434_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__nand2_1
XANTENNA__12290__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09223_ _03199_ _03229_ _04136_ _04141_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__a31o_1
X_06435_ final_design.VGA_data_control.VGA_request_address\[0\] vssd1 vssd1 vccd1
+ vccd1 _01390_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout327_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ net498 net483 vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__nor2_1
X_14220__1289 vssd1 vssd1 vccd1 vccd1 _14220__1289/HI net1289 sky130_fd_sc_hd__conb_1
XANTENNA__06653__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12952__Q net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08105_ final_design.cpu.reg_window\[972\] final_design.cpu.reg_window\[1004\] net848
+ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12593__B2 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ _02435_ net633 _04005_ net259 vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1236_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08153__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08036_ final_design.cpu.reg_window\[595\] final_design.cpu.reg_window\[627\] net825
+ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__mux2_1
Xinput90 memory_size[2] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_2
Xhold830 final_design.cpu.reg_window\[1002\] vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 final_design.cpu.reg_window\[871\] vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold852 final_design.cpu.reg_window\[395\] vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08549__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold863 final_design.cpu.reg_window\[326\] vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12390__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10356__B1 _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold874 final_design.cpu.reg_window\[795\] vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 final_design.cpu.reg_window\[429\] vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 final_design.cpu.reg_window\[129\] vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09987_ _04654_ _04656_ _04905_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout863_A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08938_ net258 _03878_ net1028 vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11305__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08869_ net632 _03815_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07524__A1 _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ net82 net1060 vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__nand2_1
XANTENNA__09712__B _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11880_ _06114_ net293 net523 net2197 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__a22o_1
XANTENNA__06828__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11871__A3 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ _05543_ _05562_ _05563_ net1018 vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13550_ clknet_leaf_117_clk _00781_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[538\]
+ sky130_fd_sc_hd__dfrtp_1
X_10762_ _05477_ _05481_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__or3_1
XANTENNA__12281__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12501_ _06163_ net354 net329 net1565 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__a22o_1
X_13481_ clknet_leaf_85_clk _00712_ net1235 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[469\]
+ sky130_fd_sc_hd__dfrtp_1
X_10693_ net977 _05432_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_62_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11322__X _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12432_ net1888 net231 net337 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__mux2_1
XANTENNA__06563__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11689__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12584__B2 final_design.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12363_ _06091_ net359 vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__and2_1
XFILLER_0_164_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ clknet_leaf_83_clk _01299_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11314_ net652 _06007_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__a21o_1
XANTENNA__09727__X _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12294_ net581 _06224_ net511 net369 net1795 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__a32o_1
XANTENNA__14171__RESET_B net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14033_ clknet_leaf_108_clk _01264_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1021\]
+ sky130_fd_sc_hd__dfrtp_1
X_11245_ _05944_ _05945_ net649 _02064_ net661 vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07394__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_X net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ final_design.reqhand.data_from_UART\[4\] net251 vssd1 vssd1 vccd1 vccd1 _05887_
+ sky130_fd_sc_hd__nand2b_2
XFILLER_0_98_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10127_ _01400_ _05000_ _05005_ vssd1 vssd1 vccd1 vccd1 final_design.v_out sky130_fd_sc_hd__or3b_1
XFILLER_0_101_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10058_ _04529_ _04530_ _04905_ _04975_ _04976_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_145_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11847__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13817_ clknet_leaf_160_clk _01048_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[805\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12272__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13748_ clknet_leaf_104_clk _00979_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[736\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10784__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13679_ clknet_leaf_94_clk _00910_ net1227 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[667\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11232__X _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11378__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07126__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08243__A2 _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07677__S1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold104 net119 vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 final_design.cpu.reg_window\[223\] vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 net126 vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09991__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold137 final_design.VGA_data_control.ready_data\[20\] vssd1 vssd1 vccd1 vccd1 net1490
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12327__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11819__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold148 final_design.cpu.reg_window\[479\] vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ net90 net93 net94 vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a21oi_1
Xhold159 final_design.reqhand.data_from_UART\[4\] vssd1 vssd1 vccd1 vccd1 net1512
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout606 net609 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_2
XANTENNA__10889__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout617 net620 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09841_ _04072_ _04753_ _04758_ _04759_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10889__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout628 net629 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_4
Xfanout639 _06157_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13894__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ net472 _04645_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06984_ _01931_ _01932_ _01933_ _01934_ net788 net794 vssd1 vssd1 vccd1 vccd1 _01935_
+ sky130_fd_sc_hd__mux4_1
X_08723_ final_design.CPU_instr_adr\[18\] _01881_ vssd1 vssd1 vccd1 vccd1 _03674_
+ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_13_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08654_ _01566_ _02604_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__nor2_1
X_07605_ _02552_ _02553_ _02554_ _02555_ net696 net715 vssd1 vssd1 vccd1 vccd1 _02556_
+ sky130_fd_sc_hd__mux4_1
X_08585_ net722 _03529_ net731 vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout444_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1186_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07536_ _02483_ _02484_ _02485_ _02486_ net780 net799 vssd1 vssd1 vccd1 vccd1 _02487_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11066__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12385__S net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07467_ _02412_ _02417_ net763 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout611_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout232_X net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09206_ _04124_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__inv_2
XFILLER_0_162_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06418_ wb_manage.curr_state\[0\] vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12015__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07398_ _02345_ _02346_ _02347_ _02348_ net785 net793 vssd1 vssd1 vccd1 vccd1 _02349_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09137_ net499 _04054_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__nand2_2
XFILLER_0_162_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1239_X net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09068_ _03786_ _03994_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12318__A1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ final_design.cpu.reg_window\[403\] final_design.cpu.reg_window\[435\] net826
+ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold660 final_design.cpu.reg_window\[470\] vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 final_design.cpu.reg_window\[427\] vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11030_ _05693_ _05709_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__nor2_1
Xhold682 final_design.cpu.reg_window\[915\] vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 final_design.cpu.reg_window\[438\] vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06412__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08103__S net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ clknet_leaf_69_clk _00212_ net1222 vssd1 vssd1 vccd1 vccd1 wb_manage.BUSY_O
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_99_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10869__A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11932_ _06133_ net282 net408 net2357 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__a22o_1
XANTENNA__10501__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ net221 net564 vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__and2_1
XFILLER_0_157_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10814_ net77 net1055 vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__nor2_1
X_13602_ clknet_leaf_23_clk _00833_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[590\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12254__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11794_ net654 net565 net200 vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__and3_1
XFILLER_0_68_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10804__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10745_ _05481_ _05482_ net1529 net1041 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_60_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13533_ clknet_leaf_32_clk _00764_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[521\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07389__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13464_ clknet_leaf_132_clk _00695_ net1167 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[452\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12006__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ net976 _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12415_ _06108_ net343 net339 net2423 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__a22o_1
X_13395_ clknet_leaf_30_clk _00626_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[383\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12346_ net2492 net360 net345 _05973_ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__a22o_1
XANTENNA__12309__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12277_ net574 _06207_ net509 net369 net1613 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__a32o_1
X_14016_ clknet_leaf_38_clk _01247_ net1136 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1004\]
+ sky130_fd_sc_hd__dfrtp_1
X_11228_ net651 _05930_ _05931_ _05932_ net662 vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__a221o_1
XANTENNA__09725__A2 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08933__B1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ final_design.reqhand.data_from_UART\[2\] net251 vssd1 vssd1 vccd1 vccd1 _05872_
+ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_147_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08948__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09633__A _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12088__A3 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11296__A1 _01881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12493__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08249__A _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11048__A1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08370_ _03308_ _03309_ _03320_ net890 vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__a22oi_4
XANTENNA__12245__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14234__1299 vssd1 vssd1 vccd1 vccd1 _14234__1299/HI net1299 sky130_fd_sc_hd__conb_1
XFILLER_0_85_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11599__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07321_ final_design.cpu.reg_window\[260\] final_design.cpu.reg_window\[292\] net940
+ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__mux2_1
XANTENNA__10032__C_N _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12260__A3 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07898__S1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06475__A1 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07252_ final_design.cpu.reg_window\[903\] final_design.cpu.reg_window\[935\] net916
+ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07672__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07183_ final_design.cpu.reg_window\[393\] final_design.cpu.reg_window\[425\] net923
+ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14022__RESET_B net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09808__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11771__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09716__A2 _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout403 _06257_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_6
Xfanout414 net415 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_8
Xfanout425 net431 vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_4
XANTENNA_fanout394_A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 _05847_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_4
X_09824_ _03262_ _04742_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__xnor2_1
Xfanout447 _04088_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_4
Xfanout458 net461 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_2
Xfanout469 net470 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07762__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10888__A1_N net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06967_ final_design.cpu.reg_window\[80\] final_design.cpu.reg_window\[112\] net958
+ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__mux2_1
X_09755_ _03229_ _04503_ _03227_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12079__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ final_design.CPU_instr_adr\[30\] _01507_ vssd1 vssd1 vccd1 vccd1 _03657_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11287__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12484__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08688__C1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09686_ net319 _04243_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__nor2_1
X_06898_ net767 _01848_ net894 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08637_ net618 _02961_ _02937_ _01938_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_7_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout826_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1189_X net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12236__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08568_ net622 net528 _03515_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__a21o_1
XANTENNA__09101__A0 final_design.CPU_instr_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07519_ _01661_ _02469_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__nor2_1
XANTENNA__07112__C1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09652__A1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08499_ _03437_ _03438_ _03449_ net892 vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12251__A3 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10530_ final_design.CPU_instr_adr\[4\] _05256_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12128__B net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10461_ net1428 net1043 _05214_ net246 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12200_ net585 _06128_ net517 net378 net2142 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__a32o_1
XANTENNA__11211__A1 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07937__S net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13180_ clknet_leaf_148_clk _00411_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[168\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_3_0_0_clk_X clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__A2 _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392_ _04991_ _05176_ _04987_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06841__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07966__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ net229 net2439 net385 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__mux2_1
XANTENNA__11459__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13745__RESET_B net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ net231 net2342 net395 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__mux2_1
Xhold490 final_design.cpu.reg_window\[787\] vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
X_11013_ _05736_ _05737_ _05719_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_53_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout970 _04043_ vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__buf_2
Xfanout981 net982 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_4
Xfanout992 _06297_ vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11278__A1 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12475__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09172__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ clknet_leaf_66_clk _00202_ net1220 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 final_design.cpu.reg_window\[164\] vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_103_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11915_ net184 _06248_ _06250_ net276 net2558 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_16_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ clknet_leaf_80_clk _00133_ net1251 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11922__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12227__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11846_ _06096_ net286 net521 net2434 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__a22o_1
XANTENNA__07329__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11777_ net2430 net412 net279 _05898_ vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__a22o_1
XFILLER_0_172_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12242__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11223__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10728_ net73 net1057 vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__nor2_1
X_13516_ clknet_leaf_118_clk _00747_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[504\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10659_ net37 _05399_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__or2_1
X_13447_ clknet_leaf_6_clk _00678_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[435\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload13 clknet_leaf_169_clk vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__inv_8
XFILLER_0_141_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload24 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__bufinv_16
Xclkload35 clknet_leaf_162_clk vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_125_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload46 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_141_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09946__A2 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ clknet_leaf_21_clk _00609_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[366\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08603__C1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload57 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload68 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_77_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload79 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_11_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12329_ net681 _05850_ _06260_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_149_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09159__B1 _01597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07148__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08057__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07870_ final_design.cpu.reg_window\[916\] final_design.cpu.reg_window\[948\] net868
+ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__mux2_1
X_06821_ final_design.cpu.reg_window\[853\] final_design.cpu.reg_window\[885\] net964
+ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__mux2_1
X_09540_ _04457_ _04458_ net477 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__mux2_1
X_06752_ net769 _01702_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__or2_1
XANTENNA__12466__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09331__B1 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09471_ _04356_ _04358_ _04388_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a21boi_1
X_06683_ final_design.cpu.reg_window\[281\] final_design.cpu.reg_window\[313\] net944
+ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11832__S net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08422_ final_design.cpu.reg_window\[837\] final_design.cpu.reg_window\[869\] net821
+ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__mux2_1
XANTENNA__12218__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09810__B _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06926__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08353_ final_design.cpu.reg_window\[7\] final_design.cpu.reg_window\[39\] net832
+ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__mux2_1
XANTENNA__06791__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12788__19 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__inv_2
XANTENNA__12229__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12233__A3 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07304_ final_design.cpu.reg_window\[837\] final_design.cpu.reg_window\[869\] net904
+ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08284_ final_design.cpu.reg_window\[457\] final_design.cpu.reg_window\[489\] net842
+ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload7 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload7/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07740__S0 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07235_ net749 _01568_ net674 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__mux2_4
XFILLER_0_61_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11992__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1149_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07166_ final_design.cpu.reg_window\[906\] final_design.cpu.reg_window\[938\] net921
+ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__mux2_1
XANTENNA__09937__A2 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07097_ final_design.cpu.reg_window\[972\] final_design.cpu.reg_window\[1004\] net929
+ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09825__X _04744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout200 _06003_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_2
Xfanout211 net212 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_2
Xfanout1209 net1217 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_2
XANTENNA_fanout776_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 _05980_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_2
Xfanout233 net234 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_2
Xfanout244 _05910_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08588__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10704__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout255 _04961_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1104_X net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09570__A0 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09273__A net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout266 net267 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_157_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09807_ net485 _04366_ _04266_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a21oi_1
Xfanout277 _06247_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_8
Xfanout288 net289 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout943_A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout299 net300 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_8
X_07999_ final_design.cpu.reg_window\[848\] final_design.cpu.reg_window\[880\] net878
+ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11308__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ net736 _04639_ _04653_ _04656_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a31o_1
XANTENNA__09858__D1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ _02801_ net441 vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11700_ net578 net422 _06208_ net296 net1755 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__a32o_1
X_12680_ _06327_ net1418 net993 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__mux2_1
XANTENNA__12209__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11631_ net210 net638 vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12224__A3 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11562_ net211 net643 vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ net979 _05261_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__or2_1
XANTENNA__11983__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13301_ clknet_leaf_28_clk _00532_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[289\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11493_ net181 net2512 net310 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13232_ clknet_leaf_115_clk _00463_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[220\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input72_A memory_size[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11697__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ _02894_ net601 vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12870__Q final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13163_ clknet_leaf_13_clk _00394_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[151\]
+ sky130_fd_sc_hd__dfrtp_1
X_10375_ net18 net1038 net1021 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1
+ vccd1 _00128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12114_ net2326 net199 net388 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13094_ clknet_leaf_170_clk _00325_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[82\]
+ sky130_fd_sc_hd__dfrtp_1
X_14233__1298 vssd1 vssd1 vccd1 vccd1 _14233__1298/HI net1298 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_72_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11917__S net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12045_ net1577 net201 net396 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09156__A3 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08498__S net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07798__S0 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09561__B1 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_161_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12879__RESET_B net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13996_ clknet_leaf_122_clk _01227_ net1197 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[984\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09313__A0 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12947_ clknet_leaf_55_clk _00185_ net1160 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12878_ clknet_leaf_79_clk _00116_ net1249 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07431__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09077__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11829_ net202 net2167 net266 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12215__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11974__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10792__A _04474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload102 clknet_leaf_123_clk vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__inv_6
XFILLER_0_153_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11240__X _05943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload113 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 clkload113/X sky130_fd_sc_hd__clkbuf_4
X_07020_ final_design.cpu.reg_window\[334\] final_design.cpu.reg_window\[366\] net934
+ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__mux2_1
XANTENNA__07577__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload124 clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 clkload124/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_153_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload135 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 clkload135/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__09919__A2 _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload146 clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 clkload146/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11187__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11726__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06602__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ final_design.CPU_instr_adr\[18\] _03793_ vssd1 vssd1 vccd1 vccd1 _03909_
+ sky130_fd_sc_hd__xnor2_2
XANTENNA__11827__S net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07922_ final_design.cpu.reg_window\[406\] final_design.cpu.reg_window\[438\] net819
+ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__mux2_1
XANTENNA__09805__B _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12687__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 final_design.cpu.reg_window\[18\] vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ _02803_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__inv_2
XANTENNA__07606__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08450__S1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ net750 net674 _01504_ _01754_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__o211a_1
X_07784_ net557 _02733_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06735_ _01668_ _01674_ _01685_ net898 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__a22oi_1
X_09523_ _04233_ _04235_ net480 vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__mux2_1
XANTENNA__12658__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_A _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1099_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ _04300_ _04303_ net476 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06666_ final_design.cpu.reg_window\[922\] final_design.cpu.reg_window\[954\] net953
+ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__mux2_1
XANTENNA__06656__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11662__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09032__S net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06764__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08405_ net536 _03354_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09385_ net539 net538 net537 net536 net457 net466 vssd1 vssd1 vccd1 vccd1 _04304_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06597_ final_design.cpu.reg_window\[348\] final_design.cpu.reg_window\[380\] net955
+ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout524_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12206__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11414__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _03274_ _03275_ _03286_ net888 vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07094__A1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11965__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08267_ final_design.cpu.reg_window\[714\] final_design.cpu.reg_window\[746\] net837
+ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__mux2_1
XANTENNA__12393__S net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_140_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_140_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1054_X net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ _02165_ _02166_ _02167_ _02168_ net778 net791 vssd1 vssd1 vccd1 vccd1 _02169_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08198_ final_design.cpu.reg_window\[782\] final_design.cpu.reg_window\[814\] net843
+ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout893_A _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07149_ _02099_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__inv_2
XANTENNA__09791__A0 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10160_ _05042_ _05054_ _05055_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[5\]
+ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 _01409_ vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__buf_2
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11737__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09138__A3 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _05000_ _05005_ _05004_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a21oi_1
Xfanout1017 _05173_ vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__buf_2
Xfanout1028 _01411_ vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1039 _05168_ vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07075__X _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__B1 _04231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06420__A final_design.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11038__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12972__RESET_B net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13850_ clknet_leaf_162_clk _01081_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[838\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10993_ net86 net1058 vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__or2_1
XANTENNA__10877__A _04598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13781_ clknet_leaf_26_clk _01012_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[769\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11472__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12732_ _06372_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12663_ final_design.VGA_data_control.ready_data\[19\] net1034 net989 final_design.data_from_mem\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11614_ net584 net423 _06164_ net301 net1540 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__a32o_1
XFILLER_0_154_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12594_ final_design.reqhand.instruction\[12\] net1011 net997 final_design.data_from_mem\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11545_ net433 net585 _06128_ net305 net1638 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_131_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07397__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11501__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11476_ net201 net2302 net307 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13215_ clknet_leaf_134_clk _00446_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[203\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10427_ _03160_ _05190_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__nor2_1
X_14195_ net1264 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XANTENNA__13007__RESET_B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10358_ net31 net1037 net1020 final_design.data_from_mem\[7\] vssd1 vssd1 vccd1 vccd1
+ _00111_ sky130_fd_sc_hd__o22a_1
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13146_ clknet_leaf_164_clk _00377_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[134\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13077_ clknet_leaf_40_clk _00308_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06691__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ net1753 net1052 vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__and2_1
XANTENNA__12669__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_125_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ net2261 net229 net397 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__mux2_1
XANTENNA__11341__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_2__f_clk_X clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06899__A1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10787__A net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13979_ clknet_leaf_155_clk _01210_ net1115 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[967\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06520_ net1051 net1008 net1005 _01470_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__o31a_1
XANTENNA__11644__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10447__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06746__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06451_ _01397_ _01400_ _01403_ _01404_ _01394_ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__a221o_2
XFILLER_0_158_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09170_ _03628_ _03650_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_118_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08121_ _02030_ net604 vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11947__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_122_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08052_ _02999_ _03000_ _03001_ _03002_ net682 net699 vssd1 vssd1 vccd1 vccd1 _03003_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_141_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07003_ net758 _01947_ net754 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__o21a_1
XANTENNA__11130__B _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06587__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08720__A final_design.CPU_instr_adr\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08954_ _03655_ _03893_ net1049 vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__o21a_1
XANTENNA__11784__C net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1014_A _05239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ _02852_ _02853_ _02854_ _02855_ net683 net699 vssd1 vssd1 vccd1 vccd1 _02856_
+ sky130_fd_sc_hd__mux4_1
X_08885_ _03773_ _03831_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout474_A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ final_design.cpu.reg_window\[789\] final_design.cpu.reg_window\[821\] net885
+ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07770__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout641_A _06157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ net728 _02717_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__or2_1
XANTENNA__12388__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09506_ _04385_ _04387_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__or2_1
X_06718_ final_design.cpu.reg_window\[344\] final_design.cpu.reg_window\[376\] net949
+ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07698_ net723 _02648_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06649_ net560 _01599_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__nand2_1
X_09437_ net735 _04333_ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__or3_2
XFILLER_0_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout906_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14232__1297 vssd1 vssd1 vccd1 vccd1 _14232__1297/HI net1297 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_23_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09368_ net86 _04193_ net87 vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_23_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11399__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11938__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ final_design.cpu.reg_window\[8\] final_design.cpu.reg_window\[40\] net838
+ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_113_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09299_ _02503_ net497 vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__nor2_2
XANTENNA_clkbuf_4_13__f_clk_X clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11330_ _04333_ _04355_ net663 vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout896_X net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11261_ net744 _03940_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09764__A0 _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10212_ final_design.uart.BAUD_counter\[4\] _05094_ net811 vssd1 vssd1 vccd1 vccd1
+ _05096_ sky130_fd_sc_hd__o21ai_1
X_13000_ net1342 _00231_ net1160 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11020__C1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11192_ final_design.reqhand.data_from_UART\[6\] net251 vssd1 vssd1 vccd1 vccd1 _05901_
+ sky130_fd_sc_hd__nand2b_2
XANTENNA__10374__B2 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11571__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ final_design.vga.h_current_state\[1\] _05011_ _05043_ vssd1 vssd1 vccd1 vccd1
+ _05044_ sky130_fd_sc_hd__or3_1
XANTENNA__06673__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A gpio_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ net677 _04991_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08414__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ clknet_leaf_113_clk _01133_ net1212 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[890\]
+ sky130_fd_sc_hd__dfrtp_1
X_13833_ clknet_leaf_88_clk _01064_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[821\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12298__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11626__A1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10400__A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13764_ clknet_leaf_98_clk _00995_ net1227 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[752\]
+ sky130_fd_sc_hd__dfrtp_1
X_10976_ _05701_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06728__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12715_ _06348_ _06352_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11215__B net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13695_ clknet_leaf_135_clk _00926_ net1167 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[683\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12646_ _06310_ net1409 net993 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11929__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_104_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12577_ net2092 _06293_ _06286_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10062__B1 _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11528_ net1686 net190 net526 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold308 final_design.cpu.reg_window\[767\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold319 final_design.cpu.reg_window\[790\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
X_14247_ net1312 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_151_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11459_ net244 net2383 net307 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12354__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ clknet_leaf_73_clk _01352_ net1244 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10365__B2 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13129_ clknet_leaf_89_clk _00360_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07156__A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 final_design.cpu.reg_window\[672\] vssd1 vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 final_design.cpu.reg_window\[102\] vssd1 vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14047__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08670_ _01481_ _01487_ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10668__A2 final_design.VGA_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09371__A _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ net613 _02570_ _02546_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07552_ net896 _02495_ _02501_ _02488_ _02489_ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__a32o_4
XANTENNA__11406__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06503_ _01375_ net1051 net1007 net1004 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__or4_2
XFILLER_0_88_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07483_ _02300_ _02433_ _02298_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__o21bai_2
XANTENNA__12290__A1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11840__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06434_ final_design.vga.h_current_state\[0\] vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
X_09222_ _04136_ _04140_ _04139_ _03133_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__a211o_1
XFILLER_0_146_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06934__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07049__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09153_ _03652_ net450 vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__nand2_4
XANTENNA__07049__B2 _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08104_ final_design.cpu.reg_window\[780\] final_design.cpu.reg_window\[812\] net847
+ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ _03785_ _04008_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08035_ final_design.cpu.reg_window\[659\] final_design.cpu.reg_window\[691\] net825
+ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__mux2_1
Xinput80 memory_size[20] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_2
XANTENNA__10980__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold820 final_design.cpu.reg_window\[670\] vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput91 memory_size[30] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08549__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 final_design.cpu.reg_window\[516\] vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 final_design.cpu.reg_window\[939\] vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07765__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09746__B1 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12345__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1229_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold853 final_design.cpu.reg_window\[259\] vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09546__A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold864 final_design.cpu.reg_window\[340\] vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 final_design.cpu.reg_window\[284\] vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10356__B2 final_design.data_from_mem\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout689_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold886 final_design.cpu.reg_window\[1017\] vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 final_design.cpu.reg_window\[496\] vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06655__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09986_ _04887_ _04904_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout1017_X net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout856_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ _02475_ _03816_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07524__A2 _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08182__C1 _01966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07819_ _02769_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__inv_2
X_08799_ _03676_ _03749_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11316__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10830_ _05543_ _05563_ _05562_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11608__B2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07005__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10761_ _05496_ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__nor2_1
XANTENNA__12281__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout909_X net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11750__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12500_ _06162_ net354 net329 net1708 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10692_ net973 _05430_ _05431_ _04042_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a22o_1
X_13480_ clknet_leaf_119_clk _00711_ net1199 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[468\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12033__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12431_ _06246_ _06260_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_134_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06416__Y _01371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12362_ net2345 net361 net349 _06090_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__a22o_1
XANTENNA__10595__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10595__B2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14101_ clknet_leaf_84_clk _01298_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11792__B1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11313_ _01823_ net649 _06005_ _06006_ net661 vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__a221o_1
XANTENNA__10890__A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12293_ net592 _06223_ net518 net371 net1720 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07675__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12336__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11244_ net752 _01480_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__nand2_2
XFILLER_0_121_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14032_ clknet_leaf_111_clk _01263_ net1211 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1020\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11175_ net747 _04016_ _05885_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a21oi_1
X_10126_ _04999_ _05033_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[8\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__10889__X _05620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08399__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ net68 _04940_ _04954_ _04956_ _04657_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__o221ai_1
XTAP_TAPCELL_ROW_69_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07704__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06723__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload0_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13816_ clknet_leaf_129_clk _01047_ net1176 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[804\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07142__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12272__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ clknet_leaf_34_clk _00978_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[735\]
+ sky130_fd_sc_hd__dfrtp_1
X_10959_ net1069 _05683_ net1013 final_design.CPU_instr_adr\[24\] vssd1 vssd1 vccd1
+ vccd1 _05687_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_46_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06754__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13678_ clknet_leaf_104_clk _00909_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[666\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12629_ final_design.VGA_data_control.ready_data\[2\] net1033 net988 final_design.data_from_mem\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07126__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11783__B1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold105 final_design.VGA_data_control.data_to_VGA\[30\] vssd1 vssd1 vccd1 vccd1 net1458
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold116 final_design.VGA_data_control.ready_data\[11\] vssd1 vssd1 vccd1 vccd1 net1469
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06885__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold127 final_design.cpu.reg_window\[221\] vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 net150 vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07585__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 net112 vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10338__B2 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09840_ _04517_ _04524_ net496 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06637__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout607 net609 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
Xfanout618 net619 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_4
Xfanout629 _02507_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08951__B2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14231__1296 vssd1 vssd1 vccd1 vccd1 _14231__1296/HI net1296 sky130_fd_sc_hd__conb_1
X_09771_ _04642_ _04644_ net477 vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__mux2_1
X_06983_ final_design.cpu.reg_window\[528\] final_design.cpu.reg_window\[560\] net958
+ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__mux2_1
XANTENNA__11835__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ final_design.CPU_instr_adr\[18\] _01881_ vssd1 vssd1 vccd1 vccd1 _03673_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08703__A1 _02510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09900__B1 _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07062__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ _02610_ _02642_ _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__and3_1
XANTENNA__10510__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10510__B2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07604_ final_design.cpu.reg_window\[157\] final_design.cpu.reg_window\[189\] net880
+ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__mux2_1
XANTENNA__11136__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08584_ net728 _03534_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10924__C_N net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07535_ final_design.cpu.reg_window\[159\] final_design.cpu.reg_window\[191\] net923
+ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12666__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1081_A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout437_A _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07466_ _02413_ _02414_ _02415_ _02416_ net786 net793 vssd1 vssd1 vccd1 vccd1 _02417_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06517__X _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06664__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06417_ net1 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09205_ _03631_ _04053_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__or2_4
XFILLER_0_107_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07397_ final_design.cpu.reg_window\[770\] final_design.cpu.reg_window\[802\] net947
+ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09967__B1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ _03629_ _04053_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__or2_2
XANTENNA__10577__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10577__B2 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12776__7 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__inv_2
X_09067_ final_design.CPU_instr_adr\[6\] _03785_ final_design.CPU_instr_adr\[7\] vssd1
+ vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09276__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08018_ final_design.cpu.reg_window\[467\] final_design.cpu.reg_window\[499\] net826
+ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__mux2_1
XANTENNA__10411__A1_N net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__A _01967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold650 final_design.cpu.reg_window\[697\] vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout973_A _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10329__B2 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 final_design.cpu.reg_window\[279\] vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold672 final_design.cpu.reg_window\[1015\] vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold683 final_design.cpu.reg_window\[419\] vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__B2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold694 final_design.cpu.reg_window\[66\] vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _03324_ net443 net439 _03326_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__o22a_1
XANTENNA__11745__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12980_ clknet_leaf_69_clk _00005_ net1221 vssd1 vssd1 vccd1 vccd1 wb_manage.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11931_ net2305 net408 _06254_ net427 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__a22o_1
XANTENNA__10501__A1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11862_ _06107_ net280 net520 net2356 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13601_ clknet_leaf_157_clk _00832_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[589\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10813_ net77 net1055 vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12254__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11793_ net2517 net412 net278 _05997_ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__a22o_1
XANTENNA__11480__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13532_ clknet_leaf_151_clk _00763_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[520\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10744_ _05478_ _05480_ net1015 vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09670__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12873__Q final_design.data_from_mem\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13463_ clknet_leaf_143_clk _00694_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[451\]
+ sky130_fd_sc_hd__dfrtp_1
X_10675_ net972 _05412_ _05415_ net968 vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__o22a_1
XFILLER_0_129_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12557__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12414_ _06243_ net500 net339 net2129 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13394_ clknet_leaf_26_clk _00625_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[382\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12345_ _06233_ net501 net361 net1863 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09186__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12276_ net579 _06206_ net511 net369 net1794 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__a32o_1
XANTENNA__08090__A _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14015_ clknet_leaf_135_clk _01246_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1003\]
+ sky130_fd_sc_hd__dfrtp_1
X_11227_ net739 _03968_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__or2_1
XANTENNA__09725__A3 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08933__A1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ net1031 net746 _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_147_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10109_ final_design.VGA_data_control.v_count\[2\] _05019_ _05022_ vssd1 vssd1 vccd1
+ vccd1 final_design.vga.v_next_count\[2\] sky130_fd_sc_hd__a21oi_1
X_11089_ final_design.CPU_instr_adr\[30\] net1014 _05807_ net1067 vssd1 vssd1 vccd1
+ vccd1 _05811_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_125_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11296__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09110__A1 final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07320_ final_design.cpu.reg_window\[324\] final_design.cpu.reg_window\[356\] net940
+ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_173_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11599__A3 _06155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09930__B1_N _04847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07251_ final_design.cpu.reg_window\[967\] final_design.cpu.reg_window\[999\] net915
+ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
XANTENNA__07672__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12548__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07182_ final_design.cpu.reg_window\[457\] final_design.cpu.reg_window\[489\] net924
+ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11756__A0 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__B net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09367__Y _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10734__S net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11220__A2 _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08204__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09716__A3 _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout404 net407 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10035__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout415 _06227_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_4
XANTENNA__08924__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout426 net431 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__buf_2
XANTENNA__09383__X _04302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _03293_ _04153_ _04154_ _03290_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__a31o_1
Xfanout437 _05847_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_4
Xfanout448 net449 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_4
Xfanout459 net460 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout387_A _06266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ _03229_ _04503_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06659__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06966_ _01913_ _01914_ _01915_ _01916_ net788 net806 vssd1 vssd1 vccd1 vccd1 _01917_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09035__S net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08705_ final_design.CPU_instr_adr\[30\] _01507_ vssd1 vssd1 vccd1 vccd1 _03656_
+ sky130_fd_sc_hd__and2_1
XANTENNA__08688__B1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09685_ net499 _04603_ _04602_ _04072_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__a211o_1
X_06897_ _01844_ _01845_ _01846_ _01847_ net775 net791 vssd1 vssd1 vccd1 vccd1 _01848_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout554_A _01750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_93_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_169_Left_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08636_ net607 _02961_ _02962_ _01938_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_90_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12236__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ net622 net528 _03515_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_7_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07518_ net557 _01690_ _02468_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08498_ _03443_ _03448_ net722 vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11995__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12997__RESET_B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07449_ _02396_ _02397_ _02398_ _02399_ net784 net802 vssd1 vssd1 vccd1 vccd1 _02400_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_135_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12539__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06871__C1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10460_ _02635_ net601 vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11747__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09119_ net978 _04037_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10391_ _05176_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__inv_2
X_12130_ _06094_ _06268_ _06267_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout976_X net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ net816 _05839_ _05841_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__and3_4
Xhold480 final_design.cpu.reg_window\[245\] vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold491 final_design.cpu.reg_window\[874\] vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ net87 net1058 vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_53_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12431__Y _06282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11328__X _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout960 net962 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_4
Xfanout971 net972 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_4
Xfanout982 _01416_ vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__buf_4
Xfanout993 _06297_ vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12868__Q final_design.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ clknet_leaf_66_clk _00201_ net1220 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_84_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold1180 final_design.cpu.reg_window\[310\] vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1191 final_design.cpu.reg_window\[876\] vssd1 vssd1 vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ final_design.cpu.reg_window\[411\] _05845_ vssd1 vssd1 vccd1 vccd1 _06250_
+ sky130_fd_sc_hd__or2_1
X_12894_ clknet_leaf_71_clk _00132_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_16_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11845_ net231 net2370 net522 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07329__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07260__Y _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11776_ net2541 net414 net288 _05891_ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__a22o_1
XANTENNA__08085__A _01785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09643__A2 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11986__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13515_ clknet_leaf_20_clk _00746_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[503\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11223__B net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10727_ net73 net1057 vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__and2_1
XANTENNA__07654__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14230__1295 vssd1 vssd1 vccd1 vccd1 _14230__1295/HI net1295 sky130_fd_sc_hd__conb_1
XFILLER_0_165_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13446_ clknet_leaf_0_clk _00677_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[434\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10658_ net37 _05399_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__nand2_1
XANTENNA__11738__A0 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload14 clknet_leaf_170_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload25 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__inv_8
XANTENNA__11202__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload36 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__08603__B1 _03524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13377_ clknet_leaf_152_clk _00608_ net1116 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[365\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09946__A3 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload47 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__clkinvlp_4
X_10589_ _05311_ _05333_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload58 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 clkload58/X sky130_fd_sc_hd__clkbuf_4
Xclkload69 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12328_ net1880 net177 net365 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12259_ net590 _06188_ net516 net374 net1555 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__a32o_1
XANTENNA__08906__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06917__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11910__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ net765 _01770_ net757 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__o21a_1
XANTENNA__13455__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06751_ _01698_ _01699_ _01700_ _01701_ net780 net799 vssd1 vssd1 vccd1 vccd1 _01702_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_75_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09331__A1 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09470_ _04356_ _04358_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__nand2_1
X_06682_ final_design.cpu.reg_window\[345\] final_design.cpu.reg_window\[377\] net944
+ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08421_ net717 _03365_ net730 vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__o21a_1
XANTENNA__12218__A1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08352_ final_design.cpu.reg_window\[71\] final_design.cpu.reg_window\[103\] net832
+ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11977__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07303_ net758 _02253_ net754 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08283_ final_design.cpu.reg_window\[265\] final_design.cpu.reg_window\[297\] net844
+ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload8 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_117_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07740__S1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07234_ net894 _02177_ _02183_ _02170_ _02171_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a32o_2
XANTENNA__06942__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07165_ final_design.cpu.reg_window\[970\] final_design.cpu.reg_window\[1002\] net921
+ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1044_A _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10401__B1 _05183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07948__A2 _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07096_ final_design.cpu.reg_window\[780\] final_design.cpu.reg_window\[812\] net928
+ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10952__A1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout201 _05996_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_2
Xfanout212 _05951_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_2
Xfanout223 net224 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_2
XANTENNA__10704__A1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 _05983_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout292_X net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout245 _05910_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_2
Xfanout256 net258 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ _04704_ _04724_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_31_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09570__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__A2 _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout267 net269 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09273__B net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 net283 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_4
X_14254__1319 vssd1 vssd1 vccd1 vccd1 _14254__1319/HI net1319 sky130_fd_sc_hd__conb_1
Xfanout289 net294 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_2
X_07998_ net723 _02942_ net731 vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__o21a_1
XANTENNA__13196__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09737_ _04184_ _04655_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__and2_1
XANTENNA__12457__A1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07008__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06949_ final_design.cpu.reg_window\[913\] final_design.cpu.reg_window\[945\] net918
+ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout936_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09668_ _04583_ _04584_ _04586_ _04342_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__o22a_1
XFILLER_0_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12209__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08619_ net542 _03194_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__nor2_1
XFILLER_0_167_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ net478 _04200_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11324__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11630_ net428 net579 _06172_ net300 net1528 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08145__A1_N net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11968__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11561_ net432 net583 _06136_ net305 net2109 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__a32o_1
XFILLER_0_92_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13300_ clknet_leaf_103_clk _00531_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[288\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10512_ final_design.CPU_instr_adr\[3\] net1014 _05255_ net1054 vssd1 vssd1 vccd1
+ vccd1 _05261_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11492_ net181 net647 vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_98_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ clknet_leaf_92_clk _00462_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[219\]
+ sky130_fd_sc_hd__dfrtp_1
X_10443_ net2460 net1047 _05205_ net248 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__a22o_1
XANTENNA__09448__B _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input65_A mem_adr_start[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ clknet_leaf_0_clk _00393_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[150\]
+ sky130_fd_sc_hd__dfrtp_1
X_10374_ net17 net1037 net1020 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1
+ vccd1 _00127_ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12113_ net1657 net201 net388 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__mux2_1
X_13093_ clknet_leaf_17_clk _00324_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07683__S net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07247__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12044_ net2044 net203 net397 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09561__A1 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07798__S1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 _01422_ vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_161_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13995_ clknet_leaf_18_clk _01226_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[983\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_57_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_161_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09313__A1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08116__A2 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12946_ clknet_leaf_56_clk _00184_ net1162 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12877_ clknet_leaf_86_clk _00115_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11234__A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11828_ net204 net2196 net266 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__mux2_1
XANTENNA__10306__S0 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11959__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11759_ net193 net2014 net417 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07858__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10792__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload103 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_116_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload114 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 clkload114/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload125 clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 clkload125/Y sky130_fd_sc_hd__clkinvlp_4
X_13429_ clknet_leaf_27_clk _00660_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[417\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload136 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 clkload136/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__11187__A1 _04863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload147 clknet_leaf_84_clk vssd1 vssd1 vccd1 vccd1 clkload147/Y sky130_fd_sc_hd__inv_6
XFILLER_0_12_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08970_ _02458_ net630 _03905_ _03907_ net256 vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__a311o_1
XANTENNA__09645__Y _04564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12136__A0 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10016__C _04934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07921_ final_design.cpu.reg_window\[470\] final_design.cpu.reg_window\[502\] net820
+ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__mux2_1
XANTENNA__13636__RESET_B net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09001__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12687__B2 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ _02800_ _02801_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__nor2_2
X_06803_ net750 net710 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__nand2_1
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
X_07783_ net621 net529 _02732_ net557 vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a211oi_1
Xclkbuf_leaf_48_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09522_ _04084_ _04440_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__and2_1
X_06734_ _01679_ _01684_ net762 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__mux2_1
XANTENNA__06937__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08718__A final_design.CPU_instr_adr\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ net492 _04342_ _04368_ _04371_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__o31a_1
X_06665_ final_design.cpu.reg_window\[986\] final_design.cpu.reg_window\[1018\] net955
+ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout252_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08404_ net619 _03352_ _03353_ _02239_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_87_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09384_ net544 net543 net541 net540 net457 net467 vssd1 vssd1 vccd1 vccd1 _04303_
+ sky130_fd_sc_hd__mux4_1
X_06596_ net771 _01546_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08335_ _03280_ _03285_ net718 vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12611__B2 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1161_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout517_A _06259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06672__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ _03213_ _03214_ _03215_ _03216_ net686 net707 vssd1 vssd1 vccd1 vccd1 _03217_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11150__Y _05864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07217_ final_design.cpu.reg_window\[8\] final_design.cpu.reg_window\[40\] net920
+ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout305_X net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ final_design.cpu.reg_window\[846\] final_design.cpu.reg_window\[878\] net843
+ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1047_X net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07148_ net542 _02098_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout886_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09791__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07079_ _01851_ _02029_ _01821_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__o21ai_4
XANTENNA__09555__Y _04474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10090_ _05004_ _05005_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__nor2_1
Xfanout1007 _01408_ vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_2
Xfanout1018 _05172_ vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_4
Xfanout1029 net1030 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09543__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11350__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11753__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06847__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13780_ clknet_leaf_106_clk _01011_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[768\]
+ sky130_fd_sc_hd__dfrtp_1
X_10992_ net86 net1059 vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__nand2_1
XANTENNA__10877__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12731_ _06368_ _06371_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_97_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12941__RESET_B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12662_ _06318_ net1433 net993 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__mux2_1
X_11613_ net240 net640 vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12602__B2 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12593_ net1417 net1009 net995 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1
+ vccd1 _01286_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11544_ net226 net644 vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12881__Q final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11475_ net202 net646 vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__and2_1
XFILLER_0_162_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13214_ clknet_leaf_22_clk _00445_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[202\]
+ sky130_fd_sc_hd__dfrtp_1
X_10426_ net1538 net1044 _05196_ net247 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_74_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input68_X net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14194_ net1263 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10916__A1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ clknet_leaf_168_clk _00376_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[133\]
+ sky130_fd_sc_hd__dfrtp_1
X_10357_ net30 net1037 net1020 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1
+ _00110_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_111_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09194__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ clknet_leaf_101_clk _00307_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08302__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _01487_ net734 _02094_ net665 vssd1 vssd1 vccd1 vccd1 final_design.cpu.Error
+ sky130_fd_sc_hd__and4_1
XANTENNA__12669__B2 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06691__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12027_ net1819 net231 net398 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__mux2_1
XANTENNA__11341__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09922__A _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07145__C _02095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13978_ clknet_leaf_160_clk _01209_ net1111 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[966\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06757__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12929_ clknet_leaf_91_clk _00167_ net1232 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_124_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06450_ final_design.vga.v_current_state\[0\] final_design.vga.v_current_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__and2b_1
XFILLER_0_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11251__X _05953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08120_ _03070_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14253__1318 vssd1 vssd1 vccd1 vccd1 _14253__1318/HI net1318 sky130_fd_sc_hd__conb_1
XFILLER_0_154_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08051_ final_design.cpu.reg_window\[274\] final_design.cpu.reg_window\[306\] net820
+ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12357__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07002_ net767 _01952_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13817__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11838__S net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06587__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08720__B _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__X _02127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _03795_ _03892_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__nor2_1
XANTENNA__10314__Y _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07904_ final_design.cpu.reg_window\[791\] final_design.cpu.reg_window\[823\] net837
+ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__mux2_1
X_08884_ _03660_ _03661_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__and2b_1
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09832__A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07835_ final_design.cpu.reg_window\[853\] final_design.cpu.reg_window\[885\] net885
+ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__mux2_1
XANTENNA__07631__S0 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout467_A _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09289__A0 _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07766_ _02713_ _02714_ _02715_ _02716_ net693 net712 vssd1 vssd1 vccd1 vccd1 _02717_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09505_ _04421_ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__xor2_1
XFILLER_0_149_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06717_ net772 _01667_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout634_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07697_ _02644_ _02645_ _02646_ _02647_ net696 net715 vssd1 vssd1 vccd1 vccd1 _02648_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09436_ net322 _04354_ _04349_ _04347_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__o211a_1
X_06648_ net752 _01598_ net672 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_136_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09367_ net738 _04280_ _04285_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__nand3_2
XANTENNA_fanout801_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06579_ final_design.cpu.reg_window\[669\] final_design.cpu.reg_window\[701\] net957
+ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__mux2_1
XANTENNA__11399__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_X net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09279__A _04177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08318_ final_design.cpu.reg_window\[72\] final_design.cpu.reg_window\[104\] net838
+ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09298_ _04119_ _04215_ _04216_ _04212_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08249_ _02128_ net604 vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12348__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ net669 _03938_ net744 vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout889_X net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10211_ _05094_ _05095_ net811 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__and3b_1
XANTENNA__08567__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11748__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11191_ net742 _04002_ _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10374__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11571__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10142_ net1063 final_design.VGA_data_control.h_count\[3\] net1062 net1061 vssd1
+ vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__o31a_1
XANTENNA__06431__A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__S net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06673__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13140__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ _01481_ net734 net253 vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__or3_1
XANTENNA__12520__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ clknet_leaf_139_clk _01132_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[889\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__X _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__A2_N _05947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ clknet_leaf_127_clk _01063_ net1193 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[820\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07262__A _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12876__Q final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13763_ clknet_leaf_6_clk _00994_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[751\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10975_ _05679_ _05681_ _05699_ _05700_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11626__A2 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10400__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12714_ final_design.VGA_data_control.v_count\[2\] _06354_ vssd1 vssd1 vccd1 vccd1
+ _06355_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_139_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06502__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11215__C net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13694_ clknet_leaf_149_clk _00925_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[682\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12645_ final_design.VGA_data_control.ready_data\[10\] net1034 net989 final_design.data_from_mem\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08805__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12576_ net1065 final_design.uart.working_data\[8\] vssd1 vssd1 vccd1 vccd1 _06293_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_124_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07201__S net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11527_ net2221 net192 net525 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12339__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14246_ net1311 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XANTENNA__13910__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold309 final_design.cpu.reg_window\[48\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11458_ net245 net646 vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13228__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ net1455 net1040 _05187_ net247 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__a22o_1
X_14177_ clknet_leaf_69_clk _01351_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11389_ net658 net180 vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__and2_1
XANTENNA__07437__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13128_ clknet_leaf_126_clk _00359_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_13059_ clknet_leaf_7_clk _00290_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[47\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1009 final_design.cpu.reg_window\[325\] vssd1 vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12511__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07443__Y _02394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ _01539_ net626 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_132_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07551_ net896 _02495_ _02501_ _02488_ _02489_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_88_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06502_ net897 _01445_ _01451_ _01439_ _01436_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__a32o_4
XFILLER_0_174_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07482_ _02332_ _02431_ _02331_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_174_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09221_ net540 _03195_ _03226_ _03197_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__o31ai_2
X_06433_ net57 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07049__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09099__A final_design.CPU_instr_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ _03645_ _03651_ net451 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10053__A1 _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08103_ final_design.cpu.reg_window\[844\] final_design.cpu.reg_window\[876\] net848
+ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10053__B2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11250__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ final_design.CPU_instr_adr\[5\] _03784_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__nor2_1
XANTENNA__10038__A _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout215_A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Left_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08034_ final_design.cpu.reg_window\[723\] final_design.cpu.reg_window\[755\] net825
+ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__mux2_1
Xinput70 memory_size[11] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09827__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput81 memory_size[21] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_130_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold810 final_design.cpu.reg_window\[405\] vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold821 final_design.cpu.reg_window\[444\] vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput92 memory_size[31] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_4
Xhold832 final_design.cpu.reg_window\[350\] vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_171_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold843 final_design.cpu.reg_window\[337\] vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09546__B _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold854 final_design.cpu.reg_window\[840\] vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10356__A2 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1124_A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 final_design.cpu.reg_window\[379\] vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 final_design.cpu.reg_window\[162\] vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07347__A _02294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11553__B2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold887 final_design.cpu.reg_window\[1019\] vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold898 final_design.cpu.reg_window\[485\] vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ net737 _04898_ _04901_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__and3_1
XANTENNA__06655__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout584_A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ _03796_ _03877_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__or2_1
XANTENNA__11305__A1 _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ _01540_ _01541_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout751_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Left_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07818_ _02766_ _02767_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_88_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08798_ _03677_ _03678_ _03747_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__nor3_1
XFILLER_0_54_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07082__A _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11608__A2 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07749_ net610 _02698_ _02674_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10760_ net42 _05483_ _05493_ _05495_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09419_ _04336_ _04337_ net474 vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10691_ _01365_ _03957_ net1070 vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_124_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11332__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12430_ net177 net646 net349 _06281_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_134_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06426__A final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10656__A1_N net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ net2426 net361 net349 _06082_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06799__A1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14100_ clknet_leaf_83_clk _01297_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ final_design.data_from_mem\[20\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06007_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07956__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12292_ net590 _06222_ net516 net370 net1769 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__a32o_1
XANTENNA__10890__B _05620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_139_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14031_ clknet_leaf_92_clk _01262_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1019\]
+ sky130_fd_sc_hd__dfrtp_1
X_11243_ net749 _01481_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ net670 _04014_ net747 vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ final_design.VGA_data_control.v_count\[8\] _05017_ _05032_ vssd1 vssd1 vccd1
+ vccd1 _05033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08399__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10056_ _04970_ _04972_ _04973_ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__or4_1
XANTENNA__11847__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output134_A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14252__1317 vssd1 vssd1 vccd1 vccd1 _14252__1317/HI net1317 sky130_fd_sc_hd__conb_1
XANTENNA__12102__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06723__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14180__RESET_B net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13815_ clknet_leaf_143_clk _01046_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[803\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13746_ clknet_leaf_39_clk _00977_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[734\]
+ sky130_fd_sc_hd__dfrtp_1
X_10958_ net978 _05685_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__nand2_1
XANTENNA__08020__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13677_ clknet_leaf_137_clk _00908_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[665\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10889_ net676 _05608_ _05619_ net977 _05618_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__o221a_2
XFILLER_0_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06582__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12628_ _06301_ net1432 net992 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12559_ _06222_ net357 net325 net2389 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold106 final_design.VGA_data_control.data_to_VGA\[7\] vssd1 vssd1 vccd1 vccd1 net1459
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold117 final_design.cpu.reg_window\[222\] vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06885__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 final_design.VGA_data_control.ready_data\[12\] vssd1 vssd1 vccd1 vccd1 net1481
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09728__A1 _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14229_ net1294 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
Xhold139 final_design.cpu.reg_window\[210\] vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06637__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout619 net620 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ _03590_ net447 _04687_ _04688_ net263 vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__o2111a_1
X_06982_ final_design.cpu.reg_window\[592\] final_design.cpu.reg_window\[624\] net958
+ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__mux2_1
X_08721_ final_design.CPU_instr_adr\[19\] _01853_ vssd1 vssd1 vccd1 vccd1 _03672_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__11299__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1190 net1191 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__clkbuf_4
X_08652_ _02706_ _03600_ _03602_ _02673_ _03601_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__a221o_1
XANTENNA__07062__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ final_design.cpu.reg_window\[221\] final_design.cpu.reg_window\[253\] net880
+ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08583_ _03530_ _03531_ _03532_ _03533_ net691 net711 vssd1 vssd1 vccd1 vccd1 _03534_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07534_ final_design.cpu.reg_window\[223\] final_design.cpu.reg_window\[255\] net923
+ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07465_ final_design.cpu.reg_window\[512\] final_design.cpu.reg_window\[544\] net951
+ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout332_A net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09204_ net488 _04077_ _04117_ _04122_ _04068_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__o311a_1
XFILLER_0_173_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06416_ net1067 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12015__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07396_ final_design.cpu.reg_window\[834\] final_design.cpu.reg_window\[866\] net947
+ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09967__A1 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09135_ _03629_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nor2_2
XANTENNA__12682__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout218_X net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11386__A1_N net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07776__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09557__A _04474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ net633 _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout799_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ final_design.cpu.reg_window\[275\] final_design.cpu.reg_window\[307\] net828
+ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 final_design.cpu.reg_window\[989\] vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold651 final_design.cpu.reg_window\[517\] vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 final_design.cpu.reg_window\[740\] vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1127_X net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold673 final_design.reqhand.instruction\[13\] vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__A2 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold684 final_design.cpu.reg_window\[691\] vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 final_design.cpu.reg_window\[913\] vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ _04180_ _04886_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__or2_1
X_08919_ _03758_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__and2_1
XANTENNA__08400__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09899_ net490 _04664_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_86_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ net565 net245 net644 vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_86_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10501__A2 _04825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout921_X net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ net430 net208 net563 net521 net1746 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__a32o_1
X_13600_ clknet_leaf_45_clk _00831_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[588\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11761__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10812_ _04452_ net251 vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06708__X _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ net2497 net412 net280 _05990_ vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ clknet_leaf_156_clk _00762_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[519\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ _05478_ _05480_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__and2_1
XFILLER_0_165_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06564__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13462_ clknet_leaf_129_clk _00693_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[450\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input95_A memory_size[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10674_ final_design.CPU_instr_adr\[11\] _03965_ net1070 vssd1 vssd1 vccd1 vccd1
+ _05415_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12006__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12413_ _06242_ net504 net342 net2348 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13393_ clknet_leaf_110_clk _00624_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[381\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09467__A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12344_ net2415 net360 net348 _05959_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12275_ net583 _06205_ net514 net370 net1766 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__a32o_1
XANTENNA__08069__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10406__A _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input50_X net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14014_ clknet_leaf_19_clk _01245_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1002\]
+ sky130_fd_sc_hd__dfrtp_1
X_11226_ net667 _03971_ net739 vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12190__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10840__S net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ net670 _04025_ net746 vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ final_design.VGA_data_control.v_count\[2\] _05019_ _05006_ vssd1 vssd1 vccd1
+ vccd1 _05022_ sky130_fd_sc_hd__o21ai_1
X_11088_ net978 _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__nand2_1
XANTENNA__11237__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ _04614_ _04615_ _04941_ _04942_ _04957_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_76_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12493__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11453__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13729_ clknet_leaf_158_clk _00960_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[717\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07250_ final_design.cpu.reg_window\[775\] final_design.cpu.reg_window\[807\] net937
+ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09949__A1 _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07181_ final_design.cpu.reg_window\[265\] final_design.cpu.reg_window\[297\] net926
+ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07596__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08281__A _02157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06632__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11508__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout405 net407 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_4
Xfanout416 net417 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__clkbuf_8
Xfanout427 net431 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_4
X_09822_ _03293_ _04153_ _04154_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__and3_1
Xfanout438 _05847_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08480__S0 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout449 net450 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_4
X_09753_ _04660_ _04661_ _04671_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08220__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06965_ final_design.cpu.reg_window\[400\] final_design.cpu.reg_window\[432\] net966
+ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout282_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ net256 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__inv_2
X_09684_ _04097_ _04205_ _04229_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06896_ final_design.cpu.reg_window\[531\] final_design.cpu.reg_window\[563\] net908
+ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__mux2_1
XANTENNA__12484__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08635_ net607 _02961_ _02962_ _01938_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__o211a_1
XANTENNA__11692__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10986__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout547_A _01937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08566_ _02394_ net614 vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_81_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12974__Q final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07360__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07517_ _01725_ _02465_ _01692_ _01724_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07112__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08497_ _03444_ _03445_ _03446_ _03447_ net692 net702 vssd1 vssd1 vccd1 vccd1 _03448_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07112__B2 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout335_X net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout714_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07448_ final_design.cpu.reg_window\[384\] final_design.cpu.reg_window\[416\] net943
+ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07379_ _01496_ net723 net679 _01484_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA_fanout502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09118_ net1068 final_design.reqhand.current_client\[1\] vssd1 vssd1 vccd1 vccd1
+ _04037_ sky130_fd_sc_hd__or2_2
XFILLER_0_72_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14251__1316 vssd1 vssd1 vccd1 vccd1 _14251__1316/HI net1316 sky130_fd_sc_hd__conb_1
X_10390_ _02028_ _03624_ _03613_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07078__Y _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09049_ _02158_ _02159_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_4__f_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_57_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12060_ net679 _05850_ _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__or3_4
Xhold470 final_design.cpu.reg_window\[214\] vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold481 final_design.cpu.reg_window\[752\] vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout969_X net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12172__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ net87 net1058 vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__and2_1
XANTENNA__11756__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold492 final_design.cpu.reg_window\[145\] vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11380__C1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout950 net956 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__clkbuf_4
Xfanout961 net962 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_2
Xfanout972 _04041_ vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__buf_4
Xfanout983 net985 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__buf_2
Xfanout994 _06297_ vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ clknet_leaf_66_clk _00200_ net1220 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09876__A0 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12475__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1170 net114 vssd1 vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1181 final_design.cpu.reg_window\[629\] vssd1 vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ net186 net2338 net277 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1192 final_design.cpu.reg_window\[825\] vssd1 vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12893_ clknet_leaf_79_clk _00131_ net1251 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11344__X _06035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11491__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ net816 _05842_ net564 vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__or3b_2
XANTENNA__12227__A2 _06155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07270__A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12884__Q final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11775_ net2458 net414 _06230_ net433 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__a22o_1
X_10726_ _05427_ _05449_ _05463_ _05447_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__o211a_1
X_13514_ clknet_leaf_2_clk _00745_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[502\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input98_X net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07654__A2 _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13445_ clknet_leaf_17_clk _00676_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[433\]
+ sky130_fd_sc_hd__dfrtp_1
X_10657_ net678 _05388_ _05398_ net979 _05397_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__o221a_1
XFILLER_0_125_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload15 clknet_leaf_171_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_140_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload26 clknet_leaf_151_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__09197__A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload37 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_106_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ clknet_leaf_27_clk _00607_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[364\]
+ sky130_fd_sc_hd__dfrtp_1
X_10588_ _05331_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06614__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload48 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload59 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__inv_6
X_12327_ net2084 net179 net365 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12258_ net593 _06187_ net518 net375 net1558 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__a32o_1
X_11209_ net745 _03987_ _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08462__S0 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12189_ net2154 net188 net382 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_166_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06917__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11910__A1 _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ final_design.cpu.reg_window\[151\] final_design.cpu.reg_window\[183\] net925
+ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__mux2_1
XANTENNA__12466__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06681_ _01627_ _01630_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__or2_1
XANTENNA__11674__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08420_ net725 _03370_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13495__RESET_B net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08351_ _03298_ _03299_ _03300_ _03301_ net685 net706 vssd1 vssd1 vccd1 vccd1 _03302_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07302_ _02249_ _02250_ _02251_ _02252_ net776 net795 vssd1 vssd1 vccd1 vccd1 _02253_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08282_ final_design.cpu.reg_window\[329\] final_design.cpu.reg_window\[361\] net843
+ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08563__X _03514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload9 clknet_leaf_164_clk vssd1 vssd1 vccd1 vccd1 clkload9/X sky130_fd_sc_hd__clkbuf_4
X_07233_ net894 _02177_ _02183_ _02170_ _02171_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a32oi_4
XANTENNA__08723__B _01881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09398__A2 _04302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07164_ final_design.cpu.reg_window\[778\] final_design.cpu.reg_window\[810\] net921
+ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10401__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07095_ final_design.cpu.reg_window\[844\] final_design.cpu.reg_window\[876\] net929
+ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08358__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09555__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 _05996_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout213 net214 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_2
Xfanout224 net225 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_2
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1204_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout246 net247 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_4
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ net736 _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__nand2_1
Xfanout257 net258 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09570__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout268 net269 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_8
Xfanout279 net283 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
X_07997_ net729 _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout664_A _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ net71 _04183_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06948_ final_design.cpu.reg_window\[977\] final_design.cpu.reg_window\[1009\] net918
+ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__mux2_1
XANTENNA__07008__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12__f_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__10468__A1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09667_ net486 _04578_ _04579_ _04585_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout831_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06879_ _01826_ _01827_ _01828_ _01829_ net775 net796 vssd1 vssd1 vccd1 vccd1 _01830_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout929_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08618_ _03426_ _03561_ _03567_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__a21o_1
XANTENNA__07884__A2 _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _04097_ _04437_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08549_ net719 _03493_ net730 vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__o21a_1
XANTENNA__11324__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ net213 net644 vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__and2_1
XANTENNA__12090__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10511_ net976 _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11491_ net182 net2438 net309 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13230_ clknet_leaf_115_clk _00461_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[218\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11340__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10442_ _02797_ net601 vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__nor2_1
XANTENNA__08125__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ clknet_leaf_95_clk _00392_ net1226 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[149\]
+ sky130_fd_sc_hd__dfrtp_1
X_10373_ net16 net1036 net1019 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1
+ vccd1 _00126_ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12112_ net2339 net203 net388 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__mux2_1
XANTENNA_input58_A mem_adr_start[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ clknet_leaf_93_clk _00323_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11339__X _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ net1537 net222 net399 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07247__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12879__Q final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout780 net781 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout791 net792 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_161_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13994_ clknet_leaf_2_clk _01225_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[982\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07552__X _02503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__A2 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11656__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10459__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ clknet_leaf_56_clk _00183_ net1162 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06758__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12110__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12876_ clknet_leaf_88_clk _00114_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_56_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09077__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11827_ net221 net2052 net269 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10306__S1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09479__X _04398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11758_ net195 net1962 net416 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__mux2_1
XANTENNA__12081__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ net71 net1057 net72 vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__or3b_1
XFILLER_0_125_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11689_ net217 net635 vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__and2_1
XANTENNA__06615__Y _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload104 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 clkload104/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12793__24 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__inv_2
Xclkload115 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload115/Y sky130_fd_sc_hd__inv_4
XTAP_TAPCELL_ROW_116_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13428_ clknet_leaf_141_clk _00659_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[416\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload126 clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 clkload126/Y sky130_fd_sc_hd__inv_6
Xclkload137 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 clkload137/Y sky130_fd_sc_hd__inv_6
Xclkload148 clknet_leaf_86_clk vssd1 vssd1 vccd1 vccd1 clkload148/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__12384__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13359_ clknet_leaf_90_clk _00590_ net1232 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[347\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07874__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09655__A _04571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07920_ final_design.cpu.reg_window\[278\] final_design.cpu.reg_window\[310\] net822
+ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__mux2_1
XANTENNA__09001__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12687__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11895__A0 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ _01784_ _02799_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__or2_1
XANTENNA__11409__B net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06802_ final_design.data_from_mem\[22\] net982 _01751_ vssd1 vssd1 vccd1 vccd1 _01753_
+ sky130_fd_sc_hd__o21ai_4
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_07782_ net610 net529 _02707_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09521_ _04201_ _04232_ net476 vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__mux2_1
X_06733_ _01680_ _01681_ _01682_ _01683_ net785 net803 vssd1 vssd1 vccd1 vccd1 _01684_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09304__A2 _03514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14250__1315 vssd1 vssd1 vccd1 vccd1 _14250__1315/HI net1315 sky130_fd_sc_hd__conb_1
XANTENNA__07315__B2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ _02768_ net440 _04369_ _02766_ _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__o221a_1
X_06664_ final_design.cpu.reg_window\[794\] final_design.cpu.reg_window\[826\] net953
+ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08403_ net608 _03352_ _03328_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09383_ net558 net556 net555 net554 net460 net470 vssd1 vssd1 vccd1 vccd1 _04302_
+ sky130_fd_sc_hd__mux4_2
X_06595_ _01542_ _01543_ _01544_ _01545_ net786 net793 vssd1 vssd1 vccd1 vccd1 _01546_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout245_A _05910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07079__B1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08334_ _03281_ _03282_ _03283_ _03284_ net698 net700 vssd1 vssd1 vccd1 vccd1 _03285_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09389__X _04308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12072__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08276__C1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06953__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08265_ final_design.cpu.reg_window\[906\] final_design.cpu.reg_window\[938\] net839
+ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout412_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1154_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07216_ final_design.cpu.reg_window\[72\] final_design.cpu.reg_window\[104\] net920
+ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08196_ net726 _03146_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12375__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07147_ _02097_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout200_X net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08043__A2 _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07078_ final_design.data_from_mem\[13\] net982 _02027_ vssd1 vssd1 vccd1 vccd1 _02029_
+ sky130_fd_sc_hd__o21ai_4
XANTENNA__09791__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout781_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout879_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10504__A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1008 _01408_ vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_1
XANTENNA__08426__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1019 net1020 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1207_X net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07003__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13346__RESET_B net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11638__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ _03070_ _04504_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__or2_1
X_10991_ _05681_ _05700_ _05716_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12730_ _06364_ _06370_ final_design.VGA_data_control.v_count\[0\] vssd1 vssd1 vccd1
+ vccd1 _06371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ final_design.VGA_data_control.ready_data\[18\] net1034 net989 final_design.data_from_mem\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11612_ net433 net585 _06163_ net301 net1466 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__a32o_1
XFILLER_0_132_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12063__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12592_ net2367 net1009 net995 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1
+ vccd1 _01285_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11543_ net434 net588 _06127_ net305 net2229 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11474_ net203 net2504 net307 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09178__C net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12366__A1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13213_ clknet_leaf_12_clk _00444_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[201\]
+ sky130_fd_sc_hd__dfrtp_1
X_10425_ _03096_ _05190_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__nor2_1
X_14193_ net1321 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_104_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10916__A2 _05620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13144_ clknet_leaf_133_clk _00375_ net1166 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[132\]
+ sky130_fd_sc_hd__dfrtp_1
X_10356_ net29 net1039 _05170_ final_design.data_from_mem\[5\] vssd1 vssd1 vccd1 vccd1
+ _00109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ clknet_leaf_33_clk _00306_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_10287_ net752 net747 _01494_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__or3_4
XANTENNA__12105__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12669__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12026_ _05839_ _06260_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__nor2_4
XANTENNA__11877__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11341__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09298__A1 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13977_ clknet_leaf_165_clk _01208_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[965\]
+ sky130_fd_sc_hd__dfrtp_1
X_12928_ clknet_leaf_98_clk _00166_ net1218 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfrtp_2
XANTENNA__07848__A2 _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12859_ clknet_leaf_79_clk _00097_ net1250 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11801__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08050_ final_design.cpu.reg_window\[338\] final_design.cpu.reg_window\[370\] net822
+ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07001_ _01948_ _01949_ _01950_ _01951_ net775 net796 vssd1 vssd1 vccd1 vccd1 _01952_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09758__C1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12363__X _06278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12109__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06587__A2 _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ final_design.CPU_instr_adr\[20\] _03794_ vssd1 vssd1 vccd1 vccd1 _03892_
+ sky130_fd_sc_hd__nor2_1
X_07903_ final_design.cpu.reg_window\[855\] final_design.cpu.reg_window\[887\] net836
+ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__mux2_1
X_08883_ final_design.CPU_instr_adr\[28\] net1029 _03827_ _03830_ vssd1 vssd1 vccd1
+ vccd1 _00239_ sky130_fd_sc_hd__a22o_1
XANTENNA__11868__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout195_A _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07834_ net729 _02778_ net732 vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06948__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07631__S1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09324__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07765_ final_design.cpu.reg_window\[152\] final_design.cpu.reg_window\[184\] net869
+ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__mux2_1
XANTENNA__09289__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_A net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09504_ _04195_ _04422_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__nand2_1
X_06716_ _01663_ _01664_ _01665_ _01666_ net785 net803 vssd1 vssd1 vccd1 vccd1 _01667_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12293__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07696_ final_design.cpu.reg_window\[411\] final_design.cpu.reg_window\[443\] net881
+ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09435_ _02900_ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__xnor2_1
X_06647_ final_design.reqhand.instruction\[27\] final_design.data_from_mem\[27\] net985
+ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__mux2_4
XANTENNA__10843__B2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout248_X net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout627_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07779__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ _04283_ _04284_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__or2_1
XANTENNA__06536__X _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06683__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06578_ final_design.cpu.reg_window\[733\] final_design.cpu.reg_window\[765\] net959
+ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08317_ _03264_ _03265_ _03266_ _03267_ net686 net706 vssd1 vssd1 vccd1 vccd1 _03268_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12596__B2 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09297_ net485 net319 _04202_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__or3_1
XANTENNA__09461__A1 _04231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1157_X net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08248_ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout996_A _06296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08179_ net604 _03129_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_132_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10210_ final_design.uart.BAUD_counter\[3\] _05093_ vssd1 vssd1 vccd1 vccd1 _05095_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_132_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11020__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11020__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ net669 _03723_ _04000_ net748 vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08972__B1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11571__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10141_ _05041_ final_design.h_out vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10072_ net986 _04038_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__or2_4
XANTENNA__11764__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ clknet_leaf_121_clk _01131_ net1197 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[888\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06858__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13831_ clknet_leaf_16_clk _01062_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[819\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10886__A1_N net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10974_ _05699_ _05700_ _05679_ _05681_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__a211oi_1
XANTENNA__11087__B2 _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12284__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13762_ clknet_leaf_23_clk _00993_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[750\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07386__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12713_ _06352_ _06353_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_139_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13693_ clknet_leaf_11_clk _00924_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[681\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11352__X _06042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12644_ _06309_ net1400 net993 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__mux2_1
XANTENNA__06593__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12892__Q final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12587__B2 final_design.data_from_mem\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12575_ net2475 _06292_ _06286_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09757__X _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11526_ net1971 net194 net524 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14245_ net1310 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
X_11457_ net237 net2372 net307 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10408_ _03384_ _05181_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__nor2_1
X_14176_ clknet_leaf_68_clk _01350_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11388_ _04324_ net665 _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08313__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10339_ net1462 net1024 net1001 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1
+ vccd1 _00096_ sky130_fd_sc_hd__a22o_1
X_13127_ clknet_leaf_7_clk _00358_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_13058_ clknet_leaf_28_clk _00289_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07518__A1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11314__A2 _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12009_ _06211_ net280 net400 net1939 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__a22o_1
XANTENNA__10431__X _05199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07550_ net769 _02500_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__or2_2
XANTENNA__12275__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06501_ net897 _01445_ _01451_ _01439_ _01436_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07481_ _02332_ _02431_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12290__A3 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07599__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09220_ _03134_ _03164_ _04137_ _04138_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__a31o_1
X_06432_ net56 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09151_ _03628_ _04053_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__or2_1
XANTENNA__09099__B net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08102_ net719 _03046_ net732 vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__o21a_1
XFILLER_0_140_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09082_ net633 _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__nor2_1
XANTENNA__11250__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08033_ net717 _02983_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__nor2_1
Xinput60 mem_adr_start[31] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_1
XFILLER_0_142_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold800 final_design.cpu.reg_window\[1016\] vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 memory_size[12] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold811 final_design.cpu.reg_window\[519\] vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput82 memory_size[22] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08731__B _02000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput93 memory_size[3] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_2
XANTENNA__11002__A1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold822 final_design.cpu.reg_window\[328\] vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11002__B2 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold833 final_design.cpu.reg_window\[263\] vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09746__A2 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08223__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold844 final_design.cpu.reg_window\[381\] vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold855 final_design.cpu.reg_window\[953\] vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 final_design.cpu.reg_window\[37\] vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__B1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11553__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold877 final_design.cpu.reg_window\[280\] vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07347__B _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13691__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold888 final_design.cpu.reg_window\[141\] vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _04902_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__inv_2
Xhold899 final_design.cpu.reg_window\[375\] vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1117_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08935_ final_design.CPU_instr_adr\[21\] _03795_ final_design.CPU_instr_adr\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11305__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout198_X net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ _03776_ _03814_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__xnor2_1
X_07817_ net558 _02765_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__or2_1
X_08797_ _03678_ _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_88_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout744_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07748_ _01630_ net621 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12266__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07679_ final_design.cpu.reg_window\[670\] final_design.cpu.reg_window\[702\] net850
+ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout911_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout532_X net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12281__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12018__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ net558 net556 net555 net554 net455 net464 vssd1 vssd1 vccd1 vccd1 _04337_
+ sky130_fd_sc_hd__mux4_1
X_10690_ _05425_ _05429_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_3__f_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09349_ _04267_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11241__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12360_ net2422 net363 net358 _06075_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11311_ net739 _03893_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__or2_1
XANTENNA__11759__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11792__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12291_ net593 _06221_ net519 net371 net1800 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__a32o_1
X_14030_ clknet_leaf_114_clk _01261_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1018\]
+ sky130_fd_sc_hd__dfrtp_1
X_11242_ net744 _03957_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11173_ net2465 net317 net423 _05884_ vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__a22o_1
XANTENNA_input40_A mem_adr_start[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ final_design.VGA_data_control.v_count\[1\] _04998_ _05031_ vssd1 vssd1 vccd1
+ vccd1 _05032_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11347__X _06038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10055_ _04701_ _04725_ _04768_ _04884_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__nand4_1
XANTENNA__12887__Q final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13814_ clknet_leaf_126_clk _01045_ net1192 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[802\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12257__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07359__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13745_ clknet_leaf_108_clk _00976_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[733\]
+ sky130_fd_sc_hd__dfrtp_1
X_10957_ _04040_ _05683_ _05684_ _04042_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08020__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12272__A3 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12009__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13676_ clknet_leaf_125_clk _00907_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[664\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_167_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10888_ net1066 _05615_ net1013 final_design.CPU_instr_adr\[21\] vssd1 vssd1 vccd1
+ vccd1 _05619_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_73_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06582__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12627_ final_design.VGA_data_control.ready_data\[1\] net1033 net988 final_design.data_from_mem\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11232__A1 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ _06221_ net359 net325 net2240 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_171_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07531__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11783__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11509_ net2181 net244 net524 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__mux2_1
X_12489_ _06149_ net355 net333 net2085 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold107 final_design.cpu.reg_window\[707\] vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold118 final_design.cpu.reg_window\[726\] vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold129 final_design.VGA_data_control.ready_data\[4\] vssd1 vssd1 vccd1 vccd1 net1482
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ net1293 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XANTENNA__13449__RESET_B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14159_ clknet_leaf_81_clk _01333_ net1248 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout609 net615 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_2
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06981_ final_design.cpu.reg_window\[656\] final_design.cpu.reg_window\[688\] net958
+ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_14__f_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ final_design.CPU_instr_adr\[19\] _01853_ vssd1 vssd1 vccd1 vccd1 _03671_
+ sky130_fd_sc_hd__or2_1
XANTENNA__12496__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1180 net1181 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_4
Xfanout1191 net1196 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__clkbuf_4
X_08651_ _01627_ _02700_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__and2_1
XANTENNA__09900__A2 _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08703__A3 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ final_design.cpu.reg_window\[29\] final_design.cpu.reg_window\[61\] net880
+ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__mux2_1
XANTENNA__12248__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08582_ final_design.cpu.reg_window\[128\] final_design.cpu.reg_window\[160\] net862
+ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__mux2_1
XANTENNA__09113__B1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07533_ final_design.cpu.reg_window\[31\] final_design.cpu.reg_window\[63\] net923
+ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XANTENNA__08467__A2 _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07464_ final_design.cpu.reg_window\[576\] final_design.cpu.reg_window\[608\] net951
+ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__mux2_1
XANTENNA__08218__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06415_ final_design.VGA_data_control.v_count\[6\] vssd1 vssd1 vccd1 vccd1 _01370_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09203_ _04106_ _04110_ _04119_ _04121_ _04115_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__o311a_1
X_07395_ final_design.cpu.reg_window\[898\] final_design.cpu.reg_window\[930\] net946
+ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10049__A _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout325_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1067_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09134_ _03647_ net666 vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_161_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12420__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09065_ _03699_ _03724_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__xor2_1
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1234_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08016_ final_design.cpu.reg_window\[339\] final_design.cpu.reg_window\[371\] net828
+ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 final_design.cpu.reg_window\[371\] vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 final_design.cpu.reg_window\[683\] vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout694_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold652 final_design.cpu.reg_window\[857\] vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 final_design.cpu.reg_window\[686\] vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold674 final_design.cpu.reg_window\[987\] vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 final_design.cpu.reg_window\[933\] vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14189__1259 vssd1 vssd1 vccd1 vccd1 _14189__1259/HI net1259 sky130_fd_sc_hd__conb_1
Xhold696 final_design.cpu.reg_window\[760\] vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07792__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09967_ net96 _04179_ net97 vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout861_A net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ _03753_ _03765_ _03761_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__a21boi_1
XANTENNA__12487__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ net477 _04814_ _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07093__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09352__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ final_design.CPU_instr_adr\[28\] final_design.CPU_instr_adr\[27\] _03799_
+ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__and3_1
XFILLER_0_169_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10501__A3 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12239__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ _06106_ net281 net520 net1955 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10811_ _05541_ _05543_ _05545_ net1041 net109 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_0_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ net2246 net415 net294 _05981_ vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06469__A1 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ clknet_leaf_160_clk _00761_ net1105 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[518\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10742_ _05458_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06437__A net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07761__S0 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06564__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10673_ net1066 _05412_ _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_153_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13461_ clknet_leaf_26_clk _00692_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[449\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07967__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12412_ _06107_ net345 net339 net2225 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__a22o_1
XANTENNA__12411__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input88_A memory_size[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ clknet_leaf_112_clk _00623_ net1212 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[380\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11489__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12343_ net2303 net361 net349 _05952_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08371__B _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12274_ net576 _06204_ net510 net368 net1697 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_79_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09186__C net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08069__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10406__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ final_design.data_from_mem\[10\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1
+ _05930_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14013_ clknet_leaf_12_clk _01244_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1001\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input43_X net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07555__X _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ net430 _05865_ net581 net315 net2254 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10107_ _05007_ _05020_ _05021_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[1\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__08727__A_N _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11518__A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11087_ net969 _05808_ _05807_ _04040_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12478__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12113__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10038_ _04954_ _04955_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_125_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11150__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_170_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12245__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11989_ _06191_ net285 net405 net1501 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13728_ clknet_leaf_37_clk _00959_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[716\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_173_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13659_ clknet_leaf_156_clk _00890_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[647\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10008__A2 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09658__A _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06781__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12402__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07180_ final_design.cpu.reg_window\[329\] final_design.cpu.reg_window\[361\] net925
+ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08281__B net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07178__A _02127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06632__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout406 net407 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__clkbuf_8
X_09821_ _03262_ _03574_ _04738_ _04739_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__a31o_1
Xfanout417 net419 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_8
Xfanout428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_4
Xfanout439 net440 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08480__S1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__C1 _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12469__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_123_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ _04072_ _04662_ _04666_ _04670_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_33_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06964_ final_design.cpu.reg_window\[464\] final_design.cpu.reg_window\[496\] net957
+ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07117__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ _02510_ _03611_ _03635_ _03653_ _03634_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__o311a_2
XANTENNA__11141__A0 final_design.reqhand.data_from_UART\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_06895_ final_design.cpu.reg_window\[595\] final_design.cpu.reg_window\[627\] net908
+ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__mux2_1
X_09683_ _03164_ _04087_ net441 _03162_ _04601_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout275_A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11692__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07912__Y _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ _03296_ _03569_ _03578_ _03584_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__a211oi_2
XANTENNA__06956__S net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_138_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _02394_ net624 vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__or2_1
XANTENNA__12236__A3 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout442_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1184_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07516_ _01725_ _02465_ _01724_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12799__30 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__inv_2
X_08496_ final_design.cpu.reg_window\[515\] final_design.cpu.reg_window\[547\] net861
+ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07112__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11995__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07447_ final_design.cpu.reg_window\[448\] final_design.cpu.reg_window\[480\] net943
+ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09839__Y _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_170_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_170_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout707_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06544__X _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07378_ final_design.reqhand.instruction\[10\] net983 _02327_ vssd1 vssd1 vccd1 vccd1
+ _02329_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09117_ net1007 net1004 net1052 vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10507__A final_design.CPU_instr_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__S net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09048_ net631 _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold460 final_design.cpu.reg_window\[231\] vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold471 final_design.cpu.reg_window\[839\] vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ _04286_ net254 _04990_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__o21a_1
Xhold482 final_design.cpu.reg_window\[606\] vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07375__X _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09573__B1 _04409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold493 final_design.cpu.reg_window\[240\] vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08411__S net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 net941 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_4
Xfanout951 net952 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_4
Xfanout962 net965 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__buf_2
Xfanout973 _04040_ vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_4
Xfanout984 net985 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_2
Xfanout995 _06296_ vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07027__S net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ clknet_leaf_57_clk _00199_ net1220 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09876__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 final_design.cpu.reg_window\[420\] vssd1 vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 final_design.cpu.reg_window\[356\] vssd1 vssd1 vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ net188 net1842 net276 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__mux2_1
Xhold1182 net158 vssd1 vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ clknet_leaf_87_clk _00130_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[26\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold1193 final_design.cpu.reg_window\[299\] vssd1 vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08647__A _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ net679 net648 vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__and2_2
XFILLER_0_157_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12227__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11073__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11435__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11774_ net656 net565 net227 vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13513_ clknet_leaf_89_clk _00744_ net1235 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[501\]
+ sky130_fd_sc_hd__dfrtp_1
X_10725_ _05425_ _05429_ _05448_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_161_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_161_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13723__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13444_ clknet_leaf_100_clk _00675_ net1188 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[432\]
+ sky130_fd_sc_hd__dfrtp_1
X_10656_ net1069 _05394_ net1014 final_design.CPU_instr_adr\[10\] vssd1 vssd1 vccd1
+ vccd1 _05398_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload16 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_8
XFILLER_0_63_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10587_ net97 final_design.VGA_adr\[5\] vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12108__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13375_ clknet_leaf_137_clk _00606_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[363\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload27 clknet_leaf_152_clk vssd1 vssd1 vccd1 vccd1 clkload27/X sky130_fd_sc_hd__clkbuf_8
Xclkload38 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__10417__A _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06929__A1_N net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload49 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_77_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12326_ net1856 net181 net367 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12257_ net589 _06186_ net516 net374 net1576 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__a32o_1
XFILLER_0_103_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09564__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ net667 _03983_ net742 vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__o21a_1
X_12188_ net1992 net190 net382 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__mux2_1
XANTENNA__08321__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11371__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08462__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11910__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11248__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ _01395_ _04037_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__nor2_1
XANTENNA__09316__A0 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09867__A1 _04125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06680_ _01627_ _01630_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__nand2_1
XANTENNA__11674__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07878__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12218__A3 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08350_ final_design.cpu.reg_window\[391\] final_design.cpu.reg_window\[423\] net834
+ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09095__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07301_ final_design.cpu.reg_window\[389\] final_design.cpu.reg_window\[421\] net906
+ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__mux2_1
XANTENNA__11977__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14188__1258 vssd1 vssd1 vccd1 vccd1 _14188__1258/HI net1258 sky130_fd_sc_hd__conb_1
X_08281_ _02157_ net619 vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_152_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_152_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11711__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07232_ net759 _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__or2_2
XFILLER_0_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06853__A1 final_design.cpu.reg_window\[820\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07400__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07163_ final_design.cpu.reg_window\[842\] final_design.cpu.reg_window\[874\] net921
+ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10401__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07094_ net761 _02038_ net755 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08358__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_2
XANTENNA__08231__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout214 _05941_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_2
XFILLER_0_100_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout392_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 _05982_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
Xfanout247 net250 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_8
X_09804_ net449 _04707_ _04717_ _04722_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__o22a_2
Xfanout258 _03654_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09570__A3 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout269 _06237_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_8
X_07996_ _02943_ _02944_ _02945_ _02946_ net696 net715 vssd1 vssd1 vccd1 vccd1 _02947_
+ sky130_fd_sc_hd__mux4_1
X_09735_ net736 _04639_ _04653_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12688__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06947_ final_design.cpu.reg_window\[785\] final_design.cpu.reg_window\[817\] net918
+ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout180_X net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09666_ net475 _04297_ net488 vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__a21oi_1
X_06878_ final_design.cpu.reg_window\[403\] final_design.cpu.reg_window\[435\] net909
+ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__mux2_1
XANTENNA__12985__Q final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08530__B2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08617_ _03426_ _03561_ _03567_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_167_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12209__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ net487 _04442_ _04515_ _04056_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1187_X net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ net727 _03498_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__or2_1
XANTENNA__11324__C net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11968__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_143_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_143_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08479_ final_design.cpu.reg_window\[387\] final_design.cpu.reg_window\[419\] net862
+ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ net971 _05255_ _05258_ net969 vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__o22a_1
X_11490_ net183 net647 vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10441_ net1444 net1048 _05204_ net248 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_98_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10928__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10372_ net15 net1038 net1021 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1
+ vccd1 _00125_ sky130_fd_sc_hd__a22o_1
X_13160_ clknet_leaf_126_clk _00391_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[148\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11767__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12111_ net1815 net222 net391 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13091_ clknet_leaf_7_clk _00322_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12042_ net2260 net205 net396 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__mux2_1
Xhold290 final_design.cpu.reg_window\[213\] vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09010__A2 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__B1 _06042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout770 _01426_ vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_2
Xfanout781 net782 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__clkbuf_8
Xfanout792 _01419_ vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__buf_8
X_13993_ clknet_leaf_85_clk _01224_ net1235 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[981\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11355__X _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12944_ clknet_leaf_56_clk _00182_ net1162 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11656__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__A3 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10459__A2 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12895__Q final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06758__S1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ clknet_leaf_86_clk _00113_ net1235 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13975__RESET_B net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11826_ net206 net2373 net266 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11959__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_134_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11757_ net196 net2334 net419 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10708_ net71 net1057 _05445_ _05446_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08316__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11688_ net427 net575 _06202_ net295 net2117 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload105 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 clkload105/X sky130_fd_sc_hd__clkbuf_8
X_13427_ clknet_leaf_31_clk _00658_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[415\]
+ sky130_fd_sc_hd__dfrtp_1
X_10639_ net814 _05378_ _05381_ _05367_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__o211a_1
Xclkload116 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 clkload116/X sky130_fd_sc_hd__clkbuf_4
Xclkload127 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 clkload127/Y sky130_fd_sc_hd__inv_6
XFILLER_0_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload138 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 clkload138/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09495__X _04414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload149 clknet_leaf_87_clk vssd1 vssd1 vccd1 vccd1 clkload149/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ clknet_leaf_113_clk _00589_ net1212 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[346\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10395__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12309_ net1978 net212 net365 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__mux2_1
XANTENNA__09655__B _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07260__B2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13289_ clknet_leaf_90_clk _00520_ net1233 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[277\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07850_ net618 _02797_ _02798_ net553 vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a211oi_2
XANTENNA__07890__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06801_ final_design.data_from_mem\[22\] net982 _01751_ vssd1 vssd1 vccd1 vccd1 _01752_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09671__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07781_ _01690_ net610 vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__and2_1
XANTENNA__06771__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_09520_ net487 _04435_ _04438_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__a21o_1
X_06732_ final_design.cpu.reg_window\[664\] final_design.cpu.reg_window\[696\] net946
+ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__mux2_1
XANTENNA__12301__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06663_ final_design.cpu.reg_window\[858\] final_design.cpu.reg_window\[890\] net953
+ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__mux2_1
X_09451_ _04085_ _04093_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07720__C1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08402_ _02240_ net621 vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06594_ final_design.cpu.reg_window\[28\] final_design.cpu.reg_window\[60\] net954
+ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__mux2_1
X_09382_ _04299_ _04300_ net476 vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08333_ final_design.cpu.reg_window\[520\] final_design.cpu.reg_window\[552\] net838
+ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__mux2_1
XANTENNA__12072__A1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_125_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08734__B _02030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout238_A _05904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ final_design.cpu.reg_window\[970\] final_design.cpu.reg_window\[1002\] net839
+ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08226__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07130__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07215_ final_design.cpu.reg_window\[136\] final_design.cpu.reg_window\[168\] net920
+ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08195_ _03142_ _03143_ _03144_ _03145_ net688 net709 vssd1 vssd1 vccd1 vccd1 _03146_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout405_A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07146_ _01503_ _02092_ _02093_ _02096_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a211o_4
XFILLER_0_14_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11583__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07077_ final_design.data_from_mem\[13\] net982 _02027_ vssd1 vssd1 vccd1 vccd1 _02028_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11277__A1_N _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09791__A3 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11159__Y _05872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1009 _06295_ vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08426__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout774_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07003__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout941_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07979_ net609 _02929_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__nor2_1
X_09718_ _04635_ _04636_ _04599_ _04616_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__a211o_1
XANTENNA__11638__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _05679_ _05700_ _05699_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_69_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09649_ _03026_ _04427_ _02996_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12660_ _06317_ net1476 net991 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11611_ net226 net640 vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12591_ net2343 net1009 net995 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1
+ vccd1 _01284_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_116_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11542_ net242 net644 vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07040__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11473_ net222 net2437 net310 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input70_A memory_size[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ clknet_leaf_147_clk _00443_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[200\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10424_ net1419 net1043 _05195_ net246 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__a22o_1
X_14192_ net1262 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_150_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10377__B2 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ clknet_leaf_144_clk _00374_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[131\]
+ sky130_fd_sc_hd__dfrtp_1
X_10355_ net28 net1037 net1020 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1
+ _00108_ sky130_fd_sc_hd__o22a_1
XANTENNA__12950__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ clknet_leaf_42_clk _00305_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_10286_ _01477_ net741 _01495_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__and3_2
XANTENNA__11326__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12025_ net816 _05841_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__nand2_4
XANTENNA__08742__A1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06753__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12121__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ clknet_leaf_131_clk _01207_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[964\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12927_ clknet_leaf_110_clk _00165_ net1214 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12858_ clknet_leaf_78_clk _00096_ net1250 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12054__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11809_ net2445 net413 net285 _06090_ vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_107_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10065__B1 _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11262__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07000_ final_design.cpu.reg_window\[143\] final_design.cpu.reg_window\[175\] net907
+ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12357__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10368__B2 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11565__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07233__A1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06667__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10605__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11200__S net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08951_ _02461_ _03889_ _03890_ net627 net256 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07902_ final_design.cpu.reg_window\[919\] final_design.cpu.reg_window\[951\] net837
+ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__mux2_1
XANTENNA__11868__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08882_ _03655_ _03829_ net1050 vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07914__A _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07092__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ net723 _02783_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08729__B _01967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout188_A _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12031__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ final_design.cpu.reg_window\[216\] final_design.cpu.reg_window\[248\] net869
+ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09503_ net88 _04194_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06715_ final_design.cpu.reg_window\[152\] final_design.cpu.reg_window\[184\] net950
+ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__mux2_1
XANTENNA__11096__A2 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12293__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07695_ final_design.cpu.reg_window\[475\] final_design.cpu.reg_window\[507\] net881
+ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout355_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09434_ _02838_ _04352_ _03036_ _03035_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06646_ net900 _01589_ _01595_ _01582_ _01583_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a32o_2
XFILLER_0_137_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09365_ _02672_ _02702_ _04282_ net450 vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout522_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06577_ net765 _01527_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_23_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08316_ final_design.cpu.reg_window\[392\] final_design.cpu.reg_window\[424\] net838
+ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09296_ _04211_ _04214_ _03485_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ _03195_ _03196_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_95_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07795__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12348__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08178_ _03116_ _03117_ _03128_ net888 vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__a22oi_4
XANTENNA__10359__B2 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout891_A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08421__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ final_design.cpu.reg_window\[843\] final_design.cpu.reg_window\[875\] net938
+ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10140_ final_design.VGA_data_control.h_count\[5\] _05014_ _05010_ final_design.vga.h_current_state\[1\]
+ final_design.vga.h_current_state\[0\] vssd1 vssd1 vccd1 vccd1 final_design.h_out
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__08972__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ net986 _04038_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11859__B2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12520__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ clknet_leaf_168_clk _01061_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[818\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13761_ clknet_leaf_158_clk _00992_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[749\]
+ sky130_fd_sc_hd__dfrtp_1
X_10973_ net84 net1059 net85 vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_67_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09685__C1 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12712_ final_design.VGA_data_control.v_count\[3\] _06351_ vssd1 vssd1 vccd1 vccd1
+ _06353_ sky130_fd_sc_hd__nand2_1
XANTENNA__07386__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08583__S0 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13692_ clknet_leaf_152_clk _00923_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[680\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08655__A _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12643_ final_design.VGA_data_control.ready_data\[9\] net1034 net989 final_design.data_from_mem\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07138__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ net1065 final_design.uart.working_data\[7\] vssd1 vssd1 vccd1 vccd1 _06292_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09452__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11525_ net2526 _06120_ _06122_ net438 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06897__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12339__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input73_X net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14244_ net1309 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11456_ net238 net646 vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__and2_1
XANTENNA__06903__A _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10407_ net1951 net1048 _05186_ net250 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14175_ clknet_leaf_68_clk _01349_ net1221 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12116__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ net660 _06070_ _06072_ _05843_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10425__A _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13126_ clknet_leaf_170_clk _00357_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_10338_ net1571 net1022 net999 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1
+ vccd1 _00095_ sky130_fd_sc_hd__a22o_1
X_13057_ clknet_leaf_159_clk _00288_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_10269_ net1626 _05129_ _05131_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12511__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07734__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ _06210_ net293 net403 net2250 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__a22o_1
XANTENNA__09912__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13237__RESET_B net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13959_ clknet_leaf_9_clk _01190_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[947\]
+ sky130_fd_sc_hd__dfrtp_1
X_06500_ net770 _01450_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07480_ _02364_ _02429_ _02362_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__o21bai_2
XANTENNA__06784__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08565__A _02394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06431_ net51 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11703__B net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09428__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09150_ _03628_ _04053_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11786__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08101_ net726 _03051_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__or2_1
X_09081_ _03705_ _03721_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__xor2_1
XANTENNA__11250__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08032_ _02979_ _02980_ _02981_ _02982_ net683 net704 vssd1 vssd1 vccd1 vccd1 _02983_
+ sky130_fd_sc_hd__mux4_1
Xinput50 mem_adr_start[22] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput61 mem_adr_start[3] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_1
Xinput72 memory_size[13] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_1
Xhold801 final_design.cpu.reg_window\[665\] vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold812 final_design.cpu.reg_window\[751\] vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 memory_size[23] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14025__RESET_B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold823 final_design.cpu.reg_window\[452\] vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput94 memory_size[4] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_2
Xhold834 final_design.cpu.reg_window\[408\] vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09600__C1 _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold845 final_design.cpu.reg_window\[523\] vssd1 vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 final_design.cpu.reg_window\[435\] vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold867 final_design.uart.BAUD_counter\[10\] vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08954__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold878 final_design.cpu.reg_window\[737\] vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ _04898_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__nand2_1
Xhold889 final_design.cpu.reg_window\[137\] vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
X_08934_ _02464_ net631 _03872_ _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1012_A _06295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07644__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ final_design.CPU_instr_adr\[29\] _01538_ vssd1 vssd1 vccd1 vccd1 _03814_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout472_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08182__A2 _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ net621 _02763_ _02764_ net558 vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a211oi_2
X_08796_ _03679_ _03740_ _03743_ _03744_ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_88_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07747_ _02685_ _02686_ _02697_ net891 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a22oi_4
XANTENNA_fanout260_X net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout737_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06694__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07678_ final_design.cpu.reg_window\[734\] final_design.cpu.reg_window\[766\] net850
+ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09417_ net561 _01566_ net560 net559 net455 net465 vssd1 vssd1 vccd1 vccd1 _04336_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__11613__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06629_ final_design.cpu.reg_window\[155\] final_design.cpu.reg_window\[187\] net960
+ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout525_X net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08317__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10029__B1 _04231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09348_ net485 net473 net530 vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11777__B1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06879__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ _04177_ _04197_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11310_ net669 _03890_ net743 vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12290_ net589 _06220_ net516 net370 net1634 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_151_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout894_X net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11241_ net669 _03955_ net744 vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_73_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12741__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ net656 net585 net226 vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10123_ final_design.VGA_data_control.v_count\[0\] final_design.VGA_data_control.v_count\[4\]
+ final_design.VGA_data_control.v_count\[2\] final_design.VGA_data_control.v_count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__and4_1
XFILLER_0_100_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10054_ net68 _04940_ _04679_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07554__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07056__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13813_ clknet_leaf_26_clk _01044_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[801\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12257__A1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11363__X _06052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07359__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13744_ clknet_leaf_115_clk _00975_ net1204 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[732\]
+ sky130_fd_sc_hd__dfrtp_1
X_10956_ _01361_ _03859_ net1071 vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07684__B2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13675_ clknet_leaf_16_clk _00906_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[663\]
+ sky130_fd_sc_hd__dfrtp_1
X_10887_ net974 _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12626_ _06300_ net1659 net991 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__mux2_1
XANTENNA__09768__X _04687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11810__Y _06237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12557_ _06220_ net356 net325 net2069 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07288__X _02239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ net1779 net238 net524 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_91_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07531__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12488_ _06148_ net345 net331 net2133 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold108 final_design.cpu.reg_window\[201\] vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ net1292 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_22_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold119 final_design.cpu.reg_window\[719\] vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11439_ net2019 net180 net314 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14158_ clknet_leaf_81_clk _01332_ net1248 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11940__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13109_ clknet_leaf_40_clk _00340_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_14089_ clknet_leaf_96_clk _01286_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_06980_ final_design.cpu.reg_window\[720\] final_design.cpu.reg_window\[752\] net958
+ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__mux2_1
XANTENNA__08149__C1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11299__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1170 net1173 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09361__A1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1181 net1189 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__clkbuf_2
X_08650_ net610 _02668_ _02643_ _01597_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__o211a_1
Xfanout1192 net1195 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__clkbuf_4
X_07601_ final_design.cpu.reg_window\[93\] final_design.cpu.reg_window\[125\] net880
+ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12248__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08581_ final_design.cpu.reg_window\[192\] final_design.cpu.reg_window\[224\] net862
+ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09113__A1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08547__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13000__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07532_ final_design.cpu.reg_window\[95\] final_design.cpu.reg_window\[127\] net923
+ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07463_ final_design.cpu.reg_window\[640\] final_design.cpu.reg_window\[672\] net951
+ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09202_ net499 net494 _04099_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__or4_1
XFILLER_0_92_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06414_ final_design.VGA_data_control.v_count\[8\] vssd1 vssd1 vccd1 vccd1 _01369_
+ sky130_fd_sc_hd__inv_2
XANTENNA__09678__X _04597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07394_ final_design.cpu.reg_window\[962\] final_design.cpu.reg_window\[994\] net946
+ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__mux2_1
XANTENNA__11759__A0 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09133_ _03607_ _04051_ _02641_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__o21a_1
XANTENNA__12420__A1 _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout220_A _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout318_A _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ _02215_ _02437_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08015_ _01853_ net606 vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold620 final_design.cpu.reg_window\[242\] vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 final_design.cpu.reg_window\[669\] vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 final_design.reqhand.instruction\[31\] vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold653 final_design.cpu.reg_window\[492\] vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 final_design.cpu.reg_window\[786\] vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07286__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold675 final_design.cpu.reg_window\[179\] vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold686 final_design.cpu.reg_window\[803\] vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold697 final_design.cpu.reg_window\[899\] vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ _04725_ _04750_ _04768_ _04884_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__and4_1
XANTENNA__06689__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1015_X net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08917_ final_design.CPU_instr_adr\[24\] net1029 _03858_ _03860_ vssd1 vssd1 vccd1
+ vccd1 _00235_ sky130_fd_sc_hd__a22o_1
X_09897_ net471 _04815_ net483 vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout854_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_96_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08848_ final_design.CPU_instr_adr\[26\] _03798_ vssd1 vssd1 vccd1 vccd1 _03799_
+ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_3_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10823__A1_N net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ _03692_ _03694_ _03729_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10810_ net1018 _05544_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__nor2_1
XANTENNA__09104__B2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ net2480 net412 net280 _05973_ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10741_ net40 _05456_ _05460_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_101_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08863__B1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07761__S1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13460_ clknet_leaf_141_clk _00691_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[448\]
+ sky130_fd_sc_hd__dfrtp_1
X_10672_ final_design.CPU_instr_adr\[11\] net1054 net814 vssd1 vssd1 vccd1 vccd1 _05413_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_153_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12411_ net207 net563 net501 net340 net2000 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10674__S net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ clknet_leaf_90_clk _00622_ net1232 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[379\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09812__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12342_ _06232_ net502 net362 net2364 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08144__S net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12273_ net577 _06203_ net512 net369 net2128 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__a32o_1
XANTENNA__13929__RESET_B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14012_ clknet_leaf_153_clk _01243_ net1118 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1000\]
+ sky130_fd_sc_hd__dfrtp_1
X_11224_ net429 net577 _05929_ net316 net1681 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__a32o_1
X_11155_ _05839_ _05866_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__nand2_4
XANTENNA__06599__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ final_design.VGA_data_control.v_count\[0\] _05017_ final_design.VGA_data_control.v_count\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__a21o_1
XANTENNA__07029__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11086_ final_design.CPU_instr_adr\[30\] _03811_ net1072 vssd1 vssd1 vccd1 vccd1
+ _05808_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_87_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10037_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__inv_2
XANTENNA__11150__A1 _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11988_ _06190_ net286 net405 net1797 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__a22o_1
XANTENNA__08319__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09646__A2 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11989__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13727_ clknet_leaf_135_clk _00958_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[715\]
+ sky130_fd_sc_hd__dfrtp_1
X_10939_ _05645_ _05662_ net243 vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__or3_1
XANTENNA__08854__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09498__X _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13658_ clknet_leaf_160_clk _00889_ net1105 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[646\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09939__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08843__A final_design.CPU_instr_adr\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12609_ net1496 net1012 net998 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1
+ vccd1 _01302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13589_ clknet_leaf_53_clk _00820_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[577\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07178__B _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10716__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11913__A0 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__B2 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout407 _06255_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_8
X_09820_ _03295_ _03569_ _03575_ net322 vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a211o_1
Xfanout418 net419 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12304__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout429 net430 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_129_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09961__X _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ net492 _04222_ _04261_ _04667_ _04669_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__o311a_1
X_06963_ final_design.cpu.reg_window\[272\] final_design.cpu.reg_window\[304\] net957
+ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_78_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_33_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08702_ _03635_ _03645_ _03650_ _03652_ net740 vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__o311a_1
XFILLER_0_146_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09682_ _03163_ net442 vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__nor2_1
XANTENNA__11141__A1 final_design.data_from_mem\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06894_ final_design.cpu.reg_window\[659\] final_design.cpu.reg_window\[691\] net908
+ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08633_ _03166_ _03581_ _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11692__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__B _02097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout268_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11444__A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07991__S1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ _02394_ net622 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_81_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07515_ _01723_ _01725_ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__nand2_1
XANTENNA__11163__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08495_ final_design.cpu.reg_window\[579\] final_design.cpu.reg_window\[611\] net861
+ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__mux2_1
XANTENNA__12641__B2 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout435_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1177_A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07446_ final_design.cpu.reg_window\[256\] final_design.cpu.reg_window\[288\] net943
+ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10347__X _05168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07377_ final_design.reqhand.instruction\[10\] net983 _02327_ vssd1 vssd1 vccd1 vccd1
+ _02328_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout602_A _05199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09116_ net1007 net1004 net1052 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10507__B net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09047_ _03728_ _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12157__A0 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold450 final_design.cpu.reg_window\[708\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout971_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11904__A0 _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 final_design.cpu.reg_window\[910\] vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold472 final_design.cpu.reg_window\[598\] vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_147_Left_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11178__X _05889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09573__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold483 final_design.cpu.reg_window\[925\] vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold494 final_design.cpu.reg_window\[138\] vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10523__A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 net932 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_4
Xfanout941 net945 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_2
Xfanout952 net956 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_4
X_09949_ _04112_ _04867_ _04443_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__o21ba_1
Xfanout963 net964 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_69_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout974 net976 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout985 net986 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__buf_2
X_12960_ clknet_leaf_57_clk _00198_ net1162 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
Xfanout996 _06296_ vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 final_design.cpu.reg_window\[97\] vssd1 vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09876__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11911_ net191 net2187 net277 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__mux2_1
Xhold1161 final_design.cpu.reg_window\[617\] vssd1 vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 final_design.cpu.reg_window\[611\] vssd1 vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12891_ clknet_leaf_79_clk _00129_ net1251 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_142_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1183 final_design.cpu.reg_window\[363\] vssd1 vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 final_design.cpu.reg_window\[52\] vssd1 vssd1 vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
X_11842_ net177 net2150 net267 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__mux2_1
XANTENNA__08139__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_156_Left_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11773_ net2447 net414 _06229_ net434 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13512_ clknet_leaf_119_clk _00743_ net1199 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[500\]
+ sky130_fd_sc_hd__dfrtp_1
X_10724_ net736 _04613_ net246 vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__and3_1
XANTENNA__06882__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13443_ clknet_leaf_2_clk _00674_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[431\]
+ sky130_fd_sc_hd__dfrtp_1
X_10655_ net979 _05396_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload17 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__clkinvlp_4
X_13374_ clknet_leaf_146_clk _00605_ net1127 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[362\]
+ sky130_fd_sc_hd__dfrtp_1
X_10586_ net97 final_design.VGA_adr\[5\] vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__nand2_1
Xclkload28 clknet_leaf_153_clk vssd1 vssd1 vccd1 vccd1 clkload28/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10417__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload39 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__clkinv_4
X_12325_ net1924 net182 net367 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_165_Left_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12256_ net584 _06185_ net503 net374 net1807 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__a32o_1
XANTENNA__06911__A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207_ _03615_ _05913_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__nor2_2
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12187_ net2157 net192 net380 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__mux2_1
XANTENNA__12124__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ _01495_ _03614_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__nor2_1
XANTENNA__07670__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09316__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _01388_ _05790_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_0_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07878__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5__f_clk_X clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06550__A1 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08049__S net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07300_ final_design.cpu.reg_window\[453\] final_design.cpu.reg_window\[485\] net905
+ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__mux2_1
X_08280_ _03195_ _03196_ _03227_ _03228_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07231_ _02178_ _02179_ _02180_ _02181_ net778 net798 vssd1 vssd1 vccd1 vccd1 _02182_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_172_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11711__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06805__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07162_ net770 _02112_ net754 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07093_ net769 _02043_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08512__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09555__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12034__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout204 _05989_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
Xfanout215 net216 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_2
Xfanout226 net227 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_2
Xfanout237 _05904_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_2
X_09803_ net322 _04721_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__nor2_1
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_4
Xfanout259 net261 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_4
X_07995_ final_design.cpu.reg_window\[144\] final_design.cpu.reg_window\[176\] net878
+ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout385_A _06266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _04124_ _04652_ _04651_ net263 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__o211ai_4
X_06946_ final_design.cpu.reg_window\[849\] final_design.cpu.reg_window\[881\] net918
+ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09858__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07652__A _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ net320 _04301_ _04305_ net321 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__a22o_1
X_06877_ final_design.cpu.reg_window\[467\] final_design.cpu.reg_window\[499\] net909
+ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout552_A _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06539__Y _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08616_ _03359_ _03564_ _03565_ _03327_ _03566_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09596_ net475 _04240_ net487 vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12614__A1 final_design.reqhand.data_from_UART\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08547_ _03494_ _03495_ _03496_ _03497_ net687 net708 vssd1 vssd1 vccd1 vccd1 _03498_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_A _02095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08478_ final_design.cpu.reg_window\[451\] final_design.cpu.reg_window\[483\] net861
+ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07429_ final_design.cpu.reg_window\[897\] final_design.cpu.reg_window\[929\] net936
+ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11621__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10440_ _02830_ net601 vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_98_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10371_ net14 net1036 net1019 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1
+ vccd1 _00124_ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ net1829 net205 net388 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09518__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13090_ clknet_leaf_30_clk _00321_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout974_X net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12041_ net1731 net208 net397 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__mux2_1
Xhold280 final_design.cpu.reg_window\[80\] vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 final_design.cpu.reg_window\[897\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11353__B2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07038__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout760 net761 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_4
Xfanout771 net773 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_4
Xfanout782 net790 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__buf_4
XANTENNA__11105__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13992_ clknet_leaf_119_clk _01223_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[980\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06877__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout793 net794 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11105__B2 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08506__C1 _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ clknet_leaf_57_clk _00181_ net1161 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11656__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08010__X _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ clknet_leaf_87_clk _00112_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11825_ net208 net2090 net267 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__mux2_1
XANTENNA__12605__B2 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10616__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11756_ net198 net2435 net419 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__mux2_1
XANTENNA__09482__A0 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12081__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10707_ net72 net1057 vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__or2_1
XFILLER_0_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12119__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ net220 net634 vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13426_ clknet_leaf_23_clk _00657_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[414\]
+ sky130_fd_sc_hd__dfrtp_1
X_10638_ net974 _05380_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload106 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 clkload106/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10147__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload117 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 clkload117/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10919__B2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload128 clknet_leaf_85_clk vssd1 vssd1 vccd1 vccd1 clkload128/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload139 clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 clkload139/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__10654__A1_N net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ clknet_leaf_139_clk _00588_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[345\]
+ sky130_fd_sc_hd__dfrtp_1
X_10569_ _05288_ _05313_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10395__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_168_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12308_ net1921 net214 net366 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08332__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13288_ clknet_leaf_119_clk _00519_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[276\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_137_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10434__Y _05201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12239_ net577 _06169_ net512 net373 net1551 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__a32o_1
XANTENNA__11344__A1 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12541__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07643__S0 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12897__RESET_B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06800_ final_design.reqhand.instruction\[22\] net983 vssd1 vssd1 vccd1 vccd1 _01751_
+ sky130_fd_sc_hd__or2_1
X_07780_ _02718_ _02719_ _02730_ net891 vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a22oi_2
XANTENNA__06787__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06771__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_06731_ final_design.cpu.reg_window\[728\] final_design.cpu.reg_window\[760\] net950
+ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__mux2_1
X_09450_ _02767_ net447 net444 vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__o21a_1
X_06662_ net763 _01606_ net756 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__o21a_1
X_08401_ net888 _03351_ _03340_ _03339_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__o2bb2a_4
X_09381_ net548 net547 net546 net545 net457 net466 vssd1 vssd1 vccd1 vccd1 _04300_
+ sky130_fd_sc_hd__mux4_1
X_06593_ final_design.cpu.reg_window\[92\] final_design.cpu.reg_window\[124\] net954
+ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08332_ final_design.cpu.reg_window\[584\] final_design.cpu.reg_window\[616\] net834
+ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__mux2_1
XANTENNA__07079__A2 _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08507__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08263_ final_design.cpu.reg_window\[778\] final_design.cpu.reg_window\[810\] net839
+ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__mux2_1
XANTENNA__11280__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12029__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07214_ final_design.cpu.reg_window\[200\] final_design.cpu.reg_window\[232\] net920
+ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12784__15 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__inv_2
XFILLER_0_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08194_ final_design.cpu.reg_window\[142\] final_design.cpu.reg_window\[174\] net844
+ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09776__A1 _04409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07145_ _01463_ _01484_ _02095_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout300_A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1042_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11583__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07076_ net1053 _01409_ _01414_ final_design.reqhand.instruction\[13\] vssd1 vssd1
+ vccd1 vccd1 _02027_ sky130_fd_sc_hd__a31o_1
XFILLER_0_113_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11169__A _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11335__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12532__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout767_A _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ net888 _02928_ _02917_ _02911_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__o2bb2a_2
X_09717_ net735 _04626_ _04630_ _04634_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__or4b_1
X_06929_ net894 _01879_ _01868_ _01862_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__11638__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout934_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__A2 _03450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09648_ _02996_ _03026_ _04427_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__and3_1
XFILLER_0_167_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _03071_ _03102_ _04496_ _03581_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_171_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11610_ net434 net588 _06162_ net301 net1765 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__a32o_1
XFILLER_0_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12590_ net1391 net1009 net995 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1
+ vccd1 _01283_ sky130_fd_sc_hd__a22o_1
XANTENNA__09464__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07321__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ net428 net581 _06126_ net304 net2075 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11472_ net205 net2471 net307 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__mux2_1
XANTENNA__13355__RESET_B net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13211_ clknet_leaf_155_clk _00442_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[199\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09767__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _03065_ _05190_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__nor2_1
X_14191_ net1261 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_151_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13142_ clknet_leaf_130_clk _00373_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[130\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input63_A mem_adr_start[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ net27 net1039 _05170_ final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1
+ _00107_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13073_ clknet_leaf_93_clk _00304_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10285_ net2552 _05139_ _05141_ net810 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__o211a_1
XANTENNA__11326__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12523__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12024_ _02295_ _05841_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_163_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12990__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08742__A2 _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09491__B _04409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08388__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06753__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 net591 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_2
X_13975_ clknet_leaf_143_clk _01206_ net1189 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[963\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12926_ clknet_leaf_11_clk _00164_ net1092 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfrtp_1
X_12857_ clknet_leaf_71_clk _00095_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11542__A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11808_ net2498 net413 net285 _06082_ vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__a22o_1
XANTENNA__08327__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07075__A1_N net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11739_ net227 net2206 net418 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11801__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09207__B1 _04125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09758__A1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ clknet_leaf_151_clk _00640_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[397\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11565__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09158__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06667__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10605__B final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ _03669_ _03752_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11317__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12514__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ final_design.cpu.reg_window\[983\] final_design.cpu.reg_window\[1015\] net836
+ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__mux2_1
X_08881_ _03800_ _03828_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11868__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07832_ _02779_ _02780_ _02781_ _02782_ net697 net716 vssd1 vssd1 vccd1 vccd1 _02783_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12312__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__B net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07092__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ final_design.cpu.reg_window\[24\] final_design.cpu.reg_window\[56\] net869
+ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__mux2_1
X_09502_ net452 _04392_ _04419_ net733 vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__a211o_2
XFILLER_0_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06714_ final_design.cpu.reg_window\[216\] final_design.cpu.reg_window\[248\] net950
+ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07694_ final_design.cpu.reg_window\[283\] final_design.cpu.reg_window\[315\] net882
+ vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07930__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ net262 _03592_ _03033_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__o21bai_2
X_06645_ net900 _01589_ _01595_ _01582_ _01583_ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__a32oi_4
XANTENNA__08745__B _02186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11452__A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ _02702_ _04282_ _02672_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08237__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06576_ _01523_ _01524_ _01525_ _01526_ net788 net806 vssd1 vssd1 vccd1 vccd1 _01527_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_111_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08315_ final_design.cpu.reg_window\[456\] final_design.cpu.reg_window\[488\] net838
+ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09997__A1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09295_ net465 _04208_ _04213_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08246_ net542 _03194_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_166_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ _03122_ _03127_ net718 vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07128_ net764 _02072_ net756 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__o21a_1
XFILLER_0_162_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08421__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07059_ final_design.cpu.reg_window\[13\] final_design.cpu.reg_window\[45\] net913
+ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__mux2_1
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_120_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12505__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ wb_manage.curr_state\[0\] net813 _04988_ _01372_ wb_manage.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11859__A2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06735__B2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11346__B net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13760_ clknet_leaf_37_clk _00991_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[748\]
+ sky130_fd_sc_hd__dfrtp_1
X_10972_ _05697_ _05698_ _05678_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08032__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12711_ final_design.VGA_data_control.v_count\[3\] _06351_ vssd1 vssd1 vccd1 vccd1
+ _06352_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13691_ clknet_leaf_155_clk _00922_ net1115 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[679\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08583__S1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12642_ _06308_ net1399 net993 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ net1873 _06291_ _06286_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11795__B2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11524_ net595 net196 _06116_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06890__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08671__A _01568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06897__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire243 _05663_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_1
XFILLER_0_108_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14243_ net1308 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
X_11455_ net223 net2300 net307 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11547__B2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ _03415_ _05181_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14174_ clknet_leaf_69_clk _01348_ net1244 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11386_ net653 _06071_ _05947_ _01538_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10425__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14181__Q final_design.VGA_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13125_ clknet_leaf_16_clk _00356_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_10337_ net1446 net1023 net1000 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1
+ vccd1 _00094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13056_ clknet_leaf_36_clk _00287_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_10268_ final_design.uart.BAUD_counter\[25\] _05129_ net809 vssd1 vssd1 vccd1 vccd1
+ _05131_ sky130_fd_sc_hd__o21ai_1
X_12007_ _06209_ net280 net400 net2374 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12132__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ _05072_ _05081_ _05084_ _05087_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__or4_1
XANTENNA__08271__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13958_ clknet_leaf_168_clk _01189_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[946\]
+ sky130_fd_sc_hd__dfrtp_1
X_12909_ clknet_leaf_10_clk _00147_ net1091 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13889_ clknet_leaf_152_clk _01120_ net1116 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[877\]
+ sky130_fd_sc_hd__dfrtp_1
X_06430_ net44 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08100_ _03047_ _03048_ _03049_ _03050_ net687 net708 vssd1 vssd1 vccd1 vccd1 _03051_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ _02270_ _02434_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08031_ final_design.cpu.reg_window\[915\] final_design.cpu.reg_window\[947\] net825
+ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput40 mem_adr_start[13] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_1
XANTENNA__06662__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07468__Y _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12307__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput51 mem_adr_start[23] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_2
Xinput62 mem_adr_start[4] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_1
Xhold802 final_design.cpu.reg_window\[415\] vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
Xinput73 memory_size[14] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_4
XANTENNA__07197__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput84 memory_size[24] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_2
Xhold813 final_design.cpu.reg_window\[946\] vssd1 vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 memory_size[5] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_2
XFILLER_0_12_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold824 final_design.cpu.reg_window\[657\] vssd1 vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold835 final_design.cpu.reg_window\[511\] vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 final_design.cpu.reg_window\[993\] vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold857 final_design.cpu.reg_window\[392\] vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08954__A2 _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09982_ _03327_ _04899_ _04900_ net449 vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__a211o_1
Xhold868 final_design.cpu.reg_window\[151\] vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 final_design.cpu.reg_window\[287\] vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08933_ net631 _03874_ _03655_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08520__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08864_ net2562 net1030 _03809_ _03813_ vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__a22o_1
XANTENNA__12042__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07815_ net611 _02763_ _02739_ net558 vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08795_ final_design.CPU_instr_adr\[16\] _01939_ vssd1 vssd1 vccd1 vccd1 _03746_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_88_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout465_A _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07746_ _02691_ _02696_ net721 vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__mux2_1
XANTENNA__12266__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07677_ _02624_ _02625_ _02626_ _02627_ net689 net710 vssd1 vssd1 vccd1 vccd1 _02628_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout632_A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06576__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ net320 _04202_ _04234_ net321 vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06628_ final_design.cpu.reg_window\[219\] final_design.cpu.reg_window\[251\] net960
+ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10029__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11226__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08317__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ net530 net485 vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06559_ _01508_ _01509_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_118_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09278_ net92 _04196_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__xor2_1
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06879__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08229_ net722 _03173_ net731 vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__o21a_1
XANTENNA__07850__C1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11529__A1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11240_ final_design.data_from_mem\[12\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1
+ _05943_ sky130_fd_sc_hd__a21o_1
XANTENNA__09874__X _04793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout887_X net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ _04825_ net665 _05843_ _05882_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_140_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10122_ _01368_ _01370_ _05027_ _05030_ _04999_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[7\]
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_98_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10053_ _04954_ _04956_ _04971_ net736 vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__a22o_1
XANTENNA__07554__B _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07056__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06708__A1 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13812_ clknet_leaf_101_clk _01043_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[800\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13717__RESET_B net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11465__A0 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07570__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10955_ _05681_ _05682_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_158_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13743_ clknet_leaf_92_clk _00974_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[731\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_158_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12009__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10886_ net973 _05615_ _05616_ net968 vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__o2bb2a_1
X_13674_ clknet_leaf_1_clk _00905_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[662\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11217__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12625_ final_design.VGA_data_control.ready_data\[0\] net1033 net987 final_design.data_from_mem\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12556_ _06219_ net354 net325 net2239 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11507_ net1839 net223 net524 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12487_ _06147_ net343 net331 net2262 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__a22o_1
XANTENNA__10436__A _03022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold109 final_design.VGA_data_control.ready_data\[24\] vssd1 vssd1 vccd1 vccd1 net1462
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14226_ net1291 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
X_11438_ net1826 net182 net313 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12193__A1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14157_ clknet_leaf_81_clk net1495 net1248 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11369_ _01599_ _05947_ _06056_ net653 vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_10_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08492__S0 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13108_ clknet_leaf_101_clk _00339_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[96\]
+ sky130_fd_sc_hd__dfrtp_1
X_14088_ clknet_leaf_96_clk _01285_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_13039_ clknet_leaf_92_clk _00270_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12496__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1160 net1163 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__buf_4
Xfanout1171 net1173 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_4
Xfanout1182 net1183 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__clkbuf_4
Xfanout1193 net1195 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__buf_2
X_07600_ _02547_ _02548_ _02549_ _02550_ net696 net703 vssd1 vssd1 vccd1 vccd1 _02551_
+ sky130_fd_sc_hd__mux4_1
X_08580_ final_design.cpu.reg_window\[0\] final_design.cpu.reg_window\[32\] net864
+ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07531_ _02478_ _02479_ _02480_ _02481_ net780 net799 vssd1 vssd1 vccd1 vccd1 _02482_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08547__S1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07462_ final_design.cpu.reg_window\[704\] final_design.cpu.reg_window\[736\] net951
+ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09201_ _03627_ _04112_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__or2_1
X_06413_ final_design.VGA_data_control.v_count\[7\] vssd1 vssd1 vccd1 vccd1 _01368_
+ sky130_fd_sc_hd__inv_2
XANTENNA__11208__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07393_ net762 _02337_ net756 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09132_ _02610_ _04050_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__and2_1
XANTENNA__08515__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12420__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09063_ final_design.CPU_instr_adr\[8\] _03990_ net1049 vssd1 vssd1 vccd1 vccd1 _00219_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12037__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout213_A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09694__X _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08014_ _01908_ _02904_ _02930_ _02964_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__o31a_1
Xhold610 final_design.cpu.reg_window\[239\] vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_163_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold621 final_design.cpu.reg_window\[283\] vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold632 final_design.cpu.reg_window\[940\] vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 final_design.cpu.reg_window\[142\] vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold654 final_design.cpu.reg_window\[360\] vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 final_design.cpu.reg_window\[261\] vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07286__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1122_A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 final_design.cpu.reg_window\[567\] vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold687 final_design.cpu.reg_window\[504\] vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11931__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07655__A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10290__S0 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold698 final_design.cpu.reg_window\[597\] vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08250__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09965_ _04788_ _04828_ _04882_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout582_A _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ net259 _03859_ net1028 vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12487__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09896_ _02126_ net539 net538 net537 net454 net463 vssd1 vssd1 vccd1 vccd1 _04815_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09352__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ final_design.CPU_instr_adr\[25\] final_design.CPU_instr_adr\[24\] _03797_
+ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_A net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06797__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08778_ _03725_ _03727_ _03695_ _03696_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__a211o_1
XANTENNA__08486__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11447__A0 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07729_ final_design.cpu.reg_window\[90\] final_design.cpu.reg_window\[122\] net872
+ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ net41 _05476_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_0_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08863__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ _05410_ _05411_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12410_ _06106_ net348 net339 net2263 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13390_ clknet_leaf_113_clk _00621_ net1212 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[378\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08076__C1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12411__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12341_ net2440 net360 net348 _05935_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__a22o_1
XANTENNA__10422__B2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12272_ net574 _06202_ net509 net369 net1877 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_79_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14011_ clknet_leaf_155_clk _01242_ net1115 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[999\]
+ sky130_fd_sc_hd__dfrtp_1
X_11223_ net655 net218 vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08160__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ _05839_ _05866_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__and2_4
XFILLER_0_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10105_ _05019_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__inv_2
X_11085_ _05801_ _05806_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07029__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12478__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ net80 _04189_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__xor2_2
XANTENNA__11686__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11150__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09726__S0 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11987_ _06189_ net293 net407 net1911 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09500__C1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13726_ clknet_leaf_19_clk _00957_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[714\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10938_ net1015 _05665_ _05666_ net1043 net2557 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__a32o_1
XANTENNA__08854__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10869_ net48 _05599_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__nor2_1
X_13657_ clknet_leaf_167_clk _00888_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[645\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11550__A net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12608_ net1412 net1009 net995 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1
+ vccd1 _01301_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08335__S net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13588_ clknet_leaf_103_clk _00819_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[576\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06644__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11610__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10413__B2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12539_ _06202_ net347 net323 net1900 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12166__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14209_ net1278 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07475__A _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08070__S net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout408 net411 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11709__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout419 _06226_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07593__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06962_ final_design.cpu.reg_window\[336\] final_design.cpu.reg_window\[368\] net957
+ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__mux2_1
X_09750_ _03198_ net446 _04222_ _04268_ _04668_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__o221a_1
XANTENNA__12469__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09690__A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ _03645_ _03651_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_33_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09681_ _03165_ _04505_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06893_ final_design.cpu.reg_window\[723\] final_design.cpu.reg_window\[755\] net908
+ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__mux2_1
XANTENNA__06779__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ net546 _03104_ _03130_ _03134_ _03582_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__o32a_1
XANTENNA__12320__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07414__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11444__B _06094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08563_ net889 _03506_ _03512_ _03499_ _03500_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__a32o_2
XANTENNA__09098__B2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07514_ _01759_ _01789_ _02463_ _01757_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_81_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11163__C net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08494_ final_design.cpu.reg_window\[643\] final_design.cpu.reg_window\[675\] net861
+ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07445_ final_design.cpu.reg_window\[320\] final_design.cpu.reg_window\[352\] net943
+ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09849__B _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1072_A final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11460__A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07376_ final_design.data_from_mem\[10\] net981 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09115_ _04034_ final_design.CPU_instr_adr\[0\] _03812_ vssd1 vssd1 vccd1 vccd1 _00209_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11601__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08073__A2 _03022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout216_X net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10507__C net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09046_ _03693_ _03695_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout797_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold440 final_design.cpu.reg_window\[349\] vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold451 final_design.cpu.reg_window\[967\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold462 final_design.cpu.reg_window\[592\] vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12999__Q final_design.CPU_instr_adr\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold473 final_design.cpu.reg_window\[92\] vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold484 final_design.cpu.reg_window\[508\] vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11619__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold495 final_design.cpu.reg_window\[759\] vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout964_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout920 net921 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_4
Xfanout931 net932 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_4
Xfanout942 net945 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_4
X_09948_ _04755_ _04866_ net487 vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__mux2_1
Xfanout953 net955 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout964 net965 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08646__A_N net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout975 net976 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout986 _01415_ vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11668__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout997 _06296_ vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__buf_2
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ net532 net459 _04061_ net468 vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 final_design.cpu.reg_window\[313\] vssd1 vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 final_design.cpu.reg_window\[113\] vssd1 vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09876__A3 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1162 final_design.cpu.reg_window\[160\] vssd1 vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ _06031_ _06248_ _06249_ net275 net2570 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__a32o_1
XANTENNA__12230__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1173 final_design.cpu.reg_window\[149\] vssd1 vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
X_12890_ clknet_leaf_87_clk _00128_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_142_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 final_design.cpu.reg_window\[661\] vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 final_design.cpu.reg_window\[558\] vssd1 vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
X_11841_ net179 net2185 net267 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ net657 net565 net242 vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__and3_1
XANTENNA__12093__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10723_ _05458_ _05459_ _05461_ net1041 net105 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__a32o_1
XFILLER_0_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13511_ clknet_leaf_6_clk _00742_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[499\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09759__B _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input93_A memory_size[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10654_ net968 _05395_ _05394_ net973 vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__a2bb2o_1
X_13442_ clknet_leaf_14_clk _00673_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[430\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13373_ clknet_leaf_14_clk _00604_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[361\]
+ sky130_fd_sc_hd__dfrtp_1
X_10585_ net737 _04903_ net249 net677 vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload18 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__bufinv_16
Xclkload29 clknet_leaf_154_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_118_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09775__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12324_ net2227 net185 net367 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12255_ net586 _06184_ net515 net374 net1554 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__a32o_1
XANTENNA__09494__B _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11206_ net249 _05854_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__nand2_1
X_12186_ net2191 net194 net380 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_166_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ final_design.CPU_instr_adr\[0\] net746 net670 _04032_ net665 vssd1 vssd1
+ vccd1 vccd1 _05852_ sky130_fd_sc_hd__a221o_1
XANTENNA__07670__S1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09316__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ net57 _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12320__A1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ _03642_ net450 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__nor2_1
XANTENNA__12140__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10331__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12084__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11831__A0 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13709_ clknet_leaf_138_clk _00940_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[697\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09669__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07230_ final_design.cpu.reg_window\[904\] final_design.cpu.reg_window\[936\] net920
+ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12387__A1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07161_ _02108_ _02109_ _02110_ _02111_ net781 net801 vssd1 vssd1 vccd1 vccd1 _02112_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07092_ _02039_ _02040_ _02041_ _02042_ net779 net800 vssd1 vssd1 vccd1 vccd1 _02043_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12315__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11347__C1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11898__A0 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08212__C1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 net206 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_2
Xfanout216 _05934_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_2
XFILLER_0_157_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout227 _05883_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_2
X_09802_ _03358_ _04720_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__xnor2_1
Xfanout238 _05904_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xfanout249 net250 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_4
X_07994_ final_design.cpu.reg_window\[208\] final_design.cpu.reg_window\[240\] net879
+ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06945_ net758 _01889_ net754 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09733_ _03071_ _04496_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout280_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout378_A net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12050__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07652__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06876_ final_design.cpu.reg_window\[275\] final_design.cpu.reg_window\[307\] net911
+ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__mux2_1
X_09664_ _04108_ _04309_ net319 vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__o21a_1
X_08615_ net537 _03297_ _03322_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__and3b_1
X_09595_ _02704_ _04049_ _04047_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08546_ final_design.cpu.reg_window\[129\] final_design.cpu.reg_window\[161\] net850
+ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__mux2_1
XANTENNA__12075__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08764__A final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11822__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08477_ final_design.cpu.reg_window\[259\] final_design.cpu.reg_window\[291\] net862
+ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout712_A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12090__A3 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07428_ final_design.cpu.reg_window\[961\] final_design.cpu.reg_window\[993\] net932
+ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10077__Y _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07359_ _02306_ _02307_ _02308_ _02309_ net784 net805 vssd1 vssd1 vccd1 vccd1 _02310_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10389__B1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10928__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ net12 net1038 net1021 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1
+ vccd1 _00123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09029_ _02445_ _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_76_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12040_ net1958 net209 net396 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__mux2_1
Xhold270 final_design.cpu.reg_window\[652\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold281 final_design.cpu.reg_window\[762\] vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11353__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 final_design.cpu.reg_window\[520\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout750 net753 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout761 net766 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13143__RESET_B net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout772 net773 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_2
X_13991_ clknet_leaf_9_clk _01222_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[979\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout783 net790 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__clkbuf_8
Xfanout794 _01419_ vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__buf_4
XFILLER_0_137_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07562__B net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09703__C1 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12942_ clknet_leaf_66_clk _00180_ net1219 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10864__A1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ clknet_leaf_73_clk _00111_ net1244 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10864__B2 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12066__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11824_ net210 net2180 net267 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__mux2_1
XANTENNA__06893__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11813__A0 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11755_ net200 net2368 net416 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__mux2_1
XANTENNA__09482__A1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12196__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10706_ net72 net1057 vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__nand2_1
XANTENNA_input96_X net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11686_ net575 net421 _06201_ net295 net1813 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__a32o_1
XFILLER_0_125_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13425_ clknet_leaf_108_clk _00656_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[413\]
+ sky130_fd_sc_hd__dfrtp_1
X_10637_ net972 _05377_ _05379_ net970 vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload107 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 clkload107/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload118 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 clkload118/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_63_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload129 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 clkload129/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_12_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10568_ _05288_ _05313_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13356_ clknet_leaf_121_clk _00587_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[344\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_168_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08993__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12307_ net1589 net216 net364 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__mux2_1
XANTENNA__12135__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10499_ net1017 _05247_ _05248_ net1045 net1422 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__a32o_1
XANTENNA__13913__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13287_ clknet_leaf_5_clk _00518_ net1096 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[275\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10444__A _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07229__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12238_ net574 _06168_ net509 net373 net1559 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__a32o_1
X_12169_ net1808 net223 net380 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__mux2_1
XANTENNA__07643__S1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06771__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06730_ final_design.cpu.reg_window\[536\] final_design.cpu.reg_window\[568\] net948
+ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06661_ net771 _01611_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__or2_1
X_08400_ _03345_ _03350_ net724 vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09380_ net553 net552 net551 net549 net457 net466 vssd1 vssd1 vccd1 vccd1 _04299_
+ sky130_fd_sc_hd__mux4_1
X_06592_ final_design.cpu.reg_window\[156\] final_design.cpu.reg_window\[188\] net954
+ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__mux2_1
XANTENNA__08584__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08331_ final_design.cpu.reg_window\[648\] final_design.cpu.reg_window\[680\] net838
+ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12072__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08262_ final_design.cpu.reg_window\[842\] final_design.cpu.reg_window\[874\] net839
+ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07213_ _02160_ _02161_ _02162_ _02163_ net782 net797 vssd1 vssd1 vccd1 vccd1 _02164_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08193_ final_design.cpu.reg_window\[206\] final_design.cpu.reg_window\[238\] net844
+ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07144_ final_design.reqhand.instruction\[7\] final_design.data_from_mem\[7\] net985
+ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__mux2_2
XFILLER_0_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06832__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07075_ net895 _02025_ _02014_ _02008_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12045__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10791__B1 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07139__S net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10073__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08759__A final_design.CPU_instr_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1202_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout662_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _02922_ _02927_ net717 vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11185__A _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ net735 _04626_ _04630_ _04633_ _04185_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__o311ai_1
X_06928_ _01873_ _01878_ net758 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__mux2_1
XANTENNA__07398__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ _04046_ _04553_ _04554_ _04564_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__a31o_1
X_06859_ final_design.cpu.reg_window\[660\] final_design.cpu.reg_window\[692\] net947
+ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout927_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09578_ _03071_ _04496_ _03580_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07602__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12599__B2 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08529_ _03474_ _03479_ net721 vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10529__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12063__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11540_ net228 net643 vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ net206 net646 vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13210_ clknet_leaf_163_clk _00441_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[198\]
+ sky130_fd_sc_hd__dfrtp_1
X_10422_ net1611 net1044 _05194_ net247 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__a22o_1
XANTENNA__12220__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14190_ net1260 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_115_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10353_ net24 net1039 _05170_ final_design.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1
+ _00106_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13141_ clknet_leaf_40_clk _00372_ net1150 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[129\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13072_ clknet_leaf_105_clk _00303_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_111_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input56_A mem_adr_start[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ final_design.uart.BAUD_counter\[31\] _05139_ vssd1 vssd1 vccd1 vccd1 _05141_
+ sky130_fd_sc_hd__nand2_1
X_12023_ _06225_ net285 net401 net2188 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_163_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08669__A _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 net581 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_4
Xfanout591 net597 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_2
XANTENNA__12287__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13974_ clknet_leaf_129_clk _01205_ net1176 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[962\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09152__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14179__Q final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ clknet_leaf_10_clk _00163_ net1092 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12856_ clknet_leaf_83_clk _00094_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11542__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11807_ net2453 net415 net293 _06075_ vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11262__A1 _02000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ net242 net2322 net418 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11669_ net817 _02358_ net815 vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__and3_4
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13408_ clknet_leaf_35_clk _00639_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[396\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12211__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07313__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11565__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13339_ clknet_leaf_153_clk _00570_ net1117 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[327\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11317__A2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07900_ net719 _02844_ net732 vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__o21a_1
XANTENNA__09682__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08880_ final_design.CPU_instr_adr\[27\] _03799_ final_design.CPU_instr_adr\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11868__A3 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07831_ final_design.cpu.reg_window\[405\] final_design.cpu.reg_window\[437\] net884
+ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__mux2_1
XANTENNA__11717__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07762_ final_design.cpu.reg_window\[88\] final_design.cpu.reg_window\[120\] net869
+ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09501_ net452 _04392_ _04419_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__a21o_1
X_06713_ final_design.cpu.reg_window\[24\] final_design.cpu.reg_window\[56\] net950
+ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__mux2_1
X_07693_ final_design.cpu.reg_window\[347\] final_design.cpu.reg_window\[379\] net882
+ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09694__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12293__A3 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06644_ net773 _01594_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__or2_1
X_09432_ _02935_ _03585_ _03589_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__or3_1
XFILLER_0_91_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11452__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09363_ _02735_ _02768_ _04281_ _02766_ _02705_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__a311o_1
X_06575_ final_design.cpu.reg_window\[925\] final_design.cpu.reg_window\[957\] net962
+ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08314_ final_design.cpu.reg_window\[264\] final_design.cpu.reg_window\[296\] net838
+ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09294_ net468 _04203_ _04207_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__or3_1
XFILLER_0_157_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_10 _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08245_ net619 _03192_ _03193_ net541 vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_62_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout410_A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06833__Y _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout508_A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12202__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ _03123_ _03124_ _03125_ _03126_ net683 net699 vssd1 vssd1 vccd1 vccd1 _03127_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09749__A2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08406__C1 _02239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08253__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10973__C_N net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07127_ net771 _02077_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10764__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07058_ final_design.cpu.reg_window\[77\] final_design.cpu.reg_window\[109\] net913
+ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__mux2_1
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XANTENNA_fanout877_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10812__A _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11627__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10971_ net85 net1059 vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__nor2_1
XANTENNA__09685__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12284__A3 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08032__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12710_ _06349_ _06350_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_67_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07696__A0 final_design.cpu.reg_window\[411\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13690_ clknet_leaf_160_clk _00921_ net1105 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[678\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06737__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_136_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ final_design.VGA_data_control.ready_data\[8\] net1034 net989 final_design.data_from_mem\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10047__A2 _04598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ final_design.uart.receiving final_design.uart.working_data\[6\] vssd1 vssd1
+ vccd1 vccd1 _06291_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_156_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08952__A final_design.CPU_instr_adr\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07543__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11795__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11523_ net2034 net197 net526 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08671__B _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14242_ net1307 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
X_11454_ net224 net646 vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__and2_1
XANTENNA__08163__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11547__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ net1677 net1048 _05185_ net250 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__a22o_1
X_14173_ clknet_leaf_72_clk _01347_ net1245 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09070__C1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11385_ final_design.data_from_mem\[29\] net236 net234 vssd1 vssd1 vccd1 vccd1 _06071_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09783__A _04697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13124_ clknet_leaf_93_clk _00355_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[112\]
+ sky130_fd_sc_hd__dfrtp_1
X_10336_ net1514 net1023 net1000 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1
+ vccd1 _00093_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11377__X _06064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ _05129_ _05130_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__nor2_1
X_13055_ clknet_leaf_133_clk _00286_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10722__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ _06208_ net284 net401 net1912 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__a22o_1
X_10198_ _05076_ _05085_ _05086_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__or3_1
XANTENNA__08271__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09007__B net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09125__B1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13957_ clknet_leaf_150_clk _01188_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[945\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12275__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12908_ clknet_leaf_10_clk _00146_ net1091 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13888_ clknet_leaf_39_clk _01119_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[876\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12839_ clknet_leaf_77_clk _00077_ net1254 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08636__C1 _01938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08862__A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11786__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08030_ final_design.cpu.reg_window\[979\] final_design.cpu.reg_window\[1011\] net825
+ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__mux2_1
XANTENNA__06662__A1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_1
XFILLER_0_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 mem_adr_start[14] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_1
XFILLER_0_4_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput52 mem_adr_start[24] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
Xinput63 mem_adr_start[5] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_1
Xhold803 final_design.cpu.reg_window\[450\] vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 memory_size[15] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_4
Xhold814 final_design.cpu.reg_window\[338\] vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput85 memory_size[25] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__buf_2
XANTENNA__09061__C1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold825 final_design.cpu.reg_window\[935\] vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08403__A2 _03352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10746__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput96 memory_size[6] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_4
Xhold836 final_design.cpu.reg_window\[500\] vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 final_design.cpu.reg_window\[1007\] vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold858 final_design.cpu.reg_window\[888\] vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09981_ _03327_ _03356_ _04706_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__and3b_1
Xhold869 final_design.cpu.reg_window\[345\] vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08932_ _03862_ _03873_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__or2_1
XANTENNA__12323__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12499__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__A2 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ _03655_ _03811_ net1050 vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o21a_1
XANTENNA__11171__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout193_A _06031_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11710__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07814_ net611 _02763_ _02739_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__o21a_1
X_08794_ _03679_ _03740_ _03743_ _03744_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_88_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07745_ _02692_ _02693_ _02694_ _02695_ net694 net703 vssd1 vssd1 vccd1 vccd1 _02696_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout360_A net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__B _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_A net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06557__A _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ final_design.cpu.reg_window\[926\] final_design.cpu.reg_window\[958\] net850
+ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07773__S0 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07152__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06576__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09415_ _04107_ _04241_ _04116_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06627_ final_design.cpu.reg_window\[27\] final_design.cpu.reg_window\[59\] net960
+ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout246_X net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout625_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11226__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06558_ _01453_ _01507_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__or2_1
XANTENNA__12423__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09346_ net473 _04075_ _04086_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__or3_1
XANTENNA__09868__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11777__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09277_ net89 net91 _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__or3_1
XFILLER_0_145_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06489_ final_design.cpu.reg_window\[862\] final_design.cpu.reg_window\[894\] net930
+ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08228_ net728 _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08159_ _03106_ _03107_ _03108_ _03109_ net683 net705 vssd1 vssd1 vccd1 vccd1 _03110_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10737__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ net660 _05879_ _05881_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ final_design.VGA_data_control.v_count\[6\] _05026_ final_design.VGA_data_control.v_count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__a21o_1
XANTENNA__12969__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10542__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07327__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ _04659_ _04676_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__nor2_1
XANTENNA__11162__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13811_ clknet_leaf_31_clk _01042_ net1139 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[799\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07851__A _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12257__A3 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11373__A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13742_ clknet_leaf_116_clk _00973_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[730\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10954_ _05676_ _05680_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_158_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13673_ clknet_leaf_94_clk _00904_ net1227 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[661\]
+ sky130_fd_sc_hd__dfrtp_1
X_10885_ final_design.CPU_instr_adr\[21\] _03887_ net1071 vssd1 vssd1 vccd1 vccd1
+ _05616_ sky130_fd_sc_hd__mux2_1
XANTENNA__13757__RESET_B net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__Y _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11217__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12624_ _05165_ net1033 vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__nor2_1
XANTENNA__09778__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12414__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12555_ _06218_ net355 net325 net2153 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11506_ net2021 net239 net526 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12486_ _06146_ net359 net334 net2340 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__a22o_1
XANTENNA__10436__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14225_ final_design.cpu.Error vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_1
X_11437_ net1904 net184 net314 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__mux2_1
XANTENNA__09594__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14156_ clknet_leaf_78_clk _01330_ net1250 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11368_ final_design.data_from_mem\[27\] net236 net234 vssd1 vssd1 vccd1 vccd1 _06056_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08492__S1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11940__A2 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13107_ clknet_leaf_33_clk _00338_ net1129 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[95\]
+ sky130_fd_sc_hd__dfrtp_1
X_10319_ net1482 net1025 net1002 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1
+ vccd1 _00076_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12143__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14087_ clknet_leaf_84_clk _01284_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10452__A _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11299_ _04451_ net659 net598 _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__o211a_4
XANTENNA__08149__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07237__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13038_ clknet_leaf_116_clk _00269_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1150 net1153 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1161 net1163 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__buf_4
Xfanout1172 net1173 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06929__X _01880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1183 net1189 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_4
Xfanout1194 net1195 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12248__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07530_ final_design.cpu.reg_window\[415\] final_design.cpu.reg_window\[447\] net923
+ vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07461_ _02408_ _02409_ _02410_ _02411_ net786 net804 vssd1 vssd1 vccd1 vccd1 _02412_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_83_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06412_ net1031 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
X_09200_ net485 _04116_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__nand2_2
XANTENNA__11208__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07392_ net772 _02342_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__or2_1
XANTENNA__12405__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09131_ _02706_ _02771_ _03594_ _03603_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__a31o_1
XANTENNA__12318__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10967__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12420__A3 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09062_ _03654_ _03987_ _03989_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_163_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08013_ _02932_ _02933_ _02963_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_114_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold600 final_design.cpu.reg_window\[489\] vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 final_design.cpu.reg_window\[998\] vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout206_A _05972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold622 final_design.cpu.reg_window\[402\] vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 final_design.cpu.reg_window\[892\] vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07936__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold644 final_design.cpu.reg_window\[849\] vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 final_design.cpu.reg_window\[180\] vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 final_design.cpu.reg_window\[93\] vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 final_design.cpu.reg_window\[646\] vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11931__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold688 final_design.cpu.reg_window\[678\] vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09964_ _04848_ _04849_ _04881_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__and3_1
XANTENNA__12053__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold699 final_design.cpu.reg_window\[336\] vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10290__S1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1115_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ final_design.CPU_instr_adr\[24\] _03797_ vssd1 vssd1 vccd1 vccd1 _03859_
+ sky130_fd_sc_hd__xnor2_1
X_09895_ _04794_ _04796_ net464 vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout196_X net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__S net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ final_design.CPU_instr_adr\[23\] _03796_ vssd1 vssd1 vccd1 vccd1 _03797_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07671__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06797__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ _03725_ _03727_ _03696_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12239__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06571__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07728_ _02675_ _02676_ _02677_ _02678_ net694 net713 vssd1 vssd1 vccd1 vccd1 _02679_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_0_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout530_X net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07659_ _02573_ _02575_ _02605_ _02607_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10670_ _05389_ _05393_ _05391_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__o21a_1
XANTENNA__13168__RESET_B net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07610__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09329_ net451 _04199_ _04245_ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__a22o_2
XFILLER_0_146_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09812__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12411__A3 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08171__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10422__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12340_ net2483 net361 net351 _05929_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_170_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12271_ net583 _06201_ net514 net368 net2279 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__a32o_1
XFILLER_0_161_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ clknet_leaf_163_clk _01241_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[998\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11222_ net598 _05926_ _05927_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__and3_2
XANTENNA__11383__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11153_ net681 _02358_ _05838_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__or3_1
X_10104_ final_design.VGA_data_control.v_count\[0\] final_design.VGA_data_control.v_count\[1\]
+ _05017_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__and3_1
X_11084_ _05804_ _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__and2b_1
XANTENNA__09879__A1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ net735 _04950_ _04952_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__or3_4
XANTENNA__11686__A1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06896__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06468__Y _01419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11986_ _06188_ net291 net406 net1721 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__a22o_1
XANTENNA__11989__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09500__B1 _04417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13725_ clknet_leaf_12_clk _00956_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[713\]
+ sky130_fd_sc_hd__dfrtp_1
X_10937_ _05643_ _05647_ _05664_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_164_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_164_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13656_ clknet_leaf_131_clk _00887_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[644\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10868_ net48 _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12607_ net1421 net1012 net998 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1
+ vccd1 _01300_ sky130_fd_sc_hd__a22o_1
XANTENNA__11550__B net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12138__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13587_ clknet_leaf_34_clk _00818_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[575\]
+ sky130_fd_sc_hd__dfrtp_1
X_10799_ _05532_ _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12538_ _06201_ net347 net324 net1977 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__a22o_1
XANTENNA__11610__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10413__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12469_ _06253_ net503 net333 net2418 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09567__A0 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14208_ net1277 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11374__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14139_ clknet_leaf_76_clk final_design.vga.h_next_count\[8\] net1253 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[8\] sky130_fd_sc_hd__dfrtp_1
Xfanout409 net411 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_4
XANTENNA__09971__A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07593__A2 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06961_ net548 _01910_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__or2_1
XANTENNA__11126__B1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08700_ _03629_ _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09680_ _04577_ _04598_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_33_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10910__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06892_ net758 _01842_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06779__S1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07976__S0 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08631_ net604 _03160_ _03135_ _01996_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__o211ai_2
XANTENNA__11725__B net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07750__C1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08562_ net889 _03506_ _03512_ _03499_ _03500_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__a32oi_2
XANTENNA__07728__S0 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07513_ _01759_ _01789_ _02463_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_81_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_155_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_155_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08493_ final_design.cpu.reg_window\[707\] final_design.cpu.reg_window\[739\] net861
+ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07444_ _02390_ _02394_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08526__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10437__A1_N net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11460__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12048__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07375_ net899 _02318_ _02324_ _02311_ _02312_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a32o_2
XFILLER_0_146_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout323_A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09114_ net629 _04032_ _04033_ _02426_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__a22o_1
XANTENNA__11601__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11887__S net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09045_ final_design.CPU_instr_adr\[10\] _03974_ net1049 vssd1 vssd1 vccd1 vccd1
+ _00221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1232_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold430 final_design.cpu.reg_window\[55\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06570__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold441 final_design.cpu.reg_window\[748\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold452 final_design.cpu.reg_window\[454\] vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11365__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout692_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11188__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 final_design.cpu.reg_window\[549\] vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 final_design.cpu.reg_window\[573\] vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1020_X net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold485 final_design.cpu.reg_window\[836\] vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11089__A2_N net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1118_X net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold496 final_design.cpu.reg_window\[330\] vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout910 net912 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_4
Xfanout921 net922 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout932 net933 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_2
X_09947_ _04710_ _04865_ net475 vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__mux2_1
Xfanout943 net944 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__clkbuf_4
Xfanout954 net955 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout957_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_X net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout965 net966 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__buf_2
Xfanout976 _04036_ vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11668__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout987 _06299_ vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_4
X_09878_ net533 net459 _04063_ net464 vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__a211o_1
Xfanout998 _06296_ vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 final_design.cpu.reg_window\[809\] vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 final_design.cpu.reg_window\[875\] vssd1 vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ final_design.CPU_instr_adr\[31\] _02504_ vssd1 vssd1 vccd1 vccd1 _03780_
+ sky130_fd_sc_hd__xnor2_1
Xhold1152 final_design.cpu.reg_window\[294\] vssd1 vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11635__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1163 final_design.cpu.reg_window\[100\] vssd1 vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1174 final_design.cpu.reg_window\[372\] vssd1 vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10340__B2 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1185 final_design.cpu.reg_window\[98\] vssd1 vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1196 final_design.CPU_instr_adr\[4\] vssd1 vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ net181 net1793 net268 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12093__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout912_X net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_146_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_146_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11771_ net2477 net413 net286 _05865_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_120_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13510_ clknet_leaf_0_clk _00741_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[498\]
+ sky130_fd_sc_hd__dfrtp_1
X_10722_ net1018 _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ clknet_leaf_151_clk _00672_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[429\]
+ sky130_fd_sc_hd__dfrtp_1
X_10653_ final_design.CPU_instr_adr\[10\] _03968_ net1071 vssd1 vssd1 vccd1 vccd1
+ _05395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input86_A memory_size[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13372_ clknet_leaf_147_clk _00603_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[360\]
+ sky130_fd_sc_hd__dfrtp_1
X_10584_ _05309_ _05327_ _05325_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_152_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08960__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload19 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_106_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12984__RESET_B net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12323_ net1768 net187 net366 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07576__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ net571 _06183_ net507 net372 net1802 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__a32o_1
XFILLER_0_32_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11205_ net248 _05854_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12185_ _06122_ net504 _06270_ net2537 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_79_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11136_ net680 _05848_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__or3_4
XANTENNA__09316__A3 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ net979 _05789_ _05787_ _05778_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__a211o_1
X_10018_ _03612_ _03635_ _04053_ _04935_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__o31a_1
XANTENNA__10331__B2 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06630__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11969_ _06171_ net288 net406 net2331 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_137_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_137_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13708_ clknet_leaf_125_clk _00939_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[696\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13639_ clknet_leaf_10_clk _00870_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[627\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11044__C1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07160_ final_design.cpu.reg_window\[138\] final_design.cpu.reg_window\[170\] net934
+ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11595__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07091_ final_design.cpu.reg_window\[140\] final_design.cpu.reg_window\[172\] net928
+ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07015__B2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout206 _05972_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
Xfanout217 net218 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
X_09801_ _03391_ _04718_ _03564_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__a21o_1
Xfanout228 net229 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_157_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout239 _05890_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_2
X_07993_ final_design.cpu.reg_window\[16\] final_design.cpu.reg_window\[48\] net879
+ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ _04117_ _04399_ _04647_ _04341_ _04650_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__o221a_2
X_06944_ net767 _01894_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09206__A _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ net497 _04581_ _04231_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a21o_1
X_06875_ final_design.cpu.reg_window\[339\] final_design.cpu.reg_window\[371\] net911
+ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__mux2_1
XANTENNA__10322__B2 final_design.data_from_mem\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout273_A _06278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08614_ net536 _03354_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__nor2_1
X_09594_ _04282_ _04512_ net450 vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08545_ final_design.cpu.reg_window\[193\] final_design.cpu.reg_window\[225\] net850
+ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__mux2_1
XANTENNA__12075__A1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_128_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1182_A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11471__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ final_design.cpu.reg_window\[323\] final_design.cpu.reg_window\[355\] net862
+ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__mux2_1
XANTENNA__08256__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07427_ final_design.cpu.reg_window\[769\] final_design.cpu.reg_window\[801\] net930
+ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout705_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07358_ final_design.cpu.reg_window\[131\] final_design.cpu.reg_window\[163\] net942
+ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10389__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07289_ net749 _01628_ net674 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__mux2_2
XFILLER_0_143_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11410__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09087__S net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09028_ _02100_ _02101_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11338__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold260 final_design.cpu.reg_window\[749\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 final_design.cpu.reg_window\[455\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 final_design.cpu.reg_window\[524\] vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold293 final_design.cpu.reg_window\[474\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12550__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09951__B1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 net742 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__clkbuf_4
Xfanout751 net753 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_1
Xfanout762 net764 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_4
XANTENNA__10550__A final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout773 _01426_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_4
X_13990_ clknet_leaf_169_clk _01221_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[978\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07335__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout784 net790 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__clkbuf_4
Xfanout795 net796 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__buf_4
X_12941_ clknet_leaf_66_clk _00179_ net1219 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10959__A1_N net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__C net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06459__B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12872_ clknet_leaf_73_clk _00110_ net1244 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_11823_ net212 net1878 net267 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__mux2_1
XANTENNA__12066__A1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11381__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11754_ net202 net2245 net416 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__mux2_1
XANTENNA__07070__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09482__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10705_ _04632_ net251 vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11685_ net245 net634 vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13424_ clknet_leaf_114_clk _00655_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[412\]
+ sky130_fd_sc_hd__dfrtp_1
X_10636_ final_design.CPU_instr_adr\[9\] _03981_ net1071 vssd1 vssd1 vccd1 vccd1 _05379_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input89_X net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08690__A _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11577__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload108 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 clkload108/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload119 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 clkload119/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13355_ clknet_leaf_21_clk _00586_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[343\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10567_ _05311_ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12306_ net2317 net218 net365 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13286_ clknet_leaf_3_clk _00517_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[274\]
+ sky130_fd_sc_hd__dfrtp_1
X_10498_ _05233_ _05246_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__nand2_1
XANTENNA__11329__B1 _06021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10444__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12237_ net583 _06167_ net514 net372 net1553 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__a32o_1
XANTENNA__10001__B1 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12541__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12168_ net2257 net239 net382 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__mux2_1
X_11119_ _05064_ _05834_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__or2_1
XANTENNA__12151__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10460__A _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12099_ net2277 net239 net391 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__mux2_1
XANTENNA__07245__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_1
XFILLER_0_160_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11843__X _06238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06660_ _01607_ _01608_ _01609_ _01610_ net786 net794 vssd1 vssd1 vccd1 vccd1 _01611_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07720__A2 _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12057__A1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06591_ final_design.cpu.reg_window\[220\] final_design.cpu.reg_window\[252\] net954
+ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08356__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08330_ final_design.cpu.reg_window\[712\] final_design.cpu.reg_window\[744\] net839
+ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08261_ net727 _03211_ net730 vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07212_ final_design.cpu.reg_window\[392\] final_design.cpu.reg_window\[424\] net920
+ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08192_ final_design.cpu.reg_window\[14\] final_design.cpu.reg_window\[46\] net844
+ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07143_ _01463_ _01484_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12326__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__C1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07074_ _02019_ _02024_ net768 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10791__B2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1028_A _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12532__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10543__A1 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout390_A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08759__B _02330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _02923_ _02924_ _02925_ _02926_ net684 net699 vssd1 vssd1 vccd1 vccd1 _02927_
+ sky130_fd_sc_hd__mux4_1
X_09715_ _04185_ _04633_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__nand2_1
X_06927_ _01874_ _01875_ _01876_ _01877_ net774 net791 vssd1 vssd1 vccd1 vccd1 _01878_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout655_A _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout276_X net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07398__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ net488 _04559_ _04560_ _04224_ _04113_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__a221o_1
X_06858_ final_design.cpu.reg_window\[724\] final_design.cpu.reg_window\[756\] net948
+ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__mux2_1
XANTENNA__06994__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12048__A1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09577_ _03231_ _04495_ _03572_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_171_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06789_ final_design.cpu.reg_window\[726\] final_design.cpu.reg_window\[758\] net902
+ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08528_ _03475_ _03476_ _03477_ _03478_ net693 net702 vssd1 vssd1 vccd1 vccd1 _03479_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11271__A2 _05967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ final_design.cpu.reg_window\[644\] final_design.cpu.reg_window\[676\] net858
+ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11470_ net207 net2394 net308 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_6__f_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11559__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ _03192_ _05190_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12220__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ clknet_leaf_102_clk _00371_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[128\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10352_ net13 net1039 _05170_ final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1
+ _00105_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08015__A _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10782__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10782__B2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13071_ clknet_leaf_92_clk _00302_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_10283_ _05139_ _05140_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__nor2_1
X_12022_ _06224_ net286 net401 net2255 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__a22o_1
XANTENNA__12523__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input49_A mem_adr_start[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10534__A1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08669__B _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07065__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 net572 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout581 net582 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__buf_2
Xfanout592 net594 vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_4
X_13973_ clknet_leaf_26_clk _01204_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[961\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12287__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ clknet_leaf_90_clk _00162_ net1233 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12039__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12855_ clknet_leaf_82_clk _00093_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11806_ net2247 net414 net291 _06068_ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11798__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11262__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11737_ net228 net2320 net416 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__mux2_1
XANTENNA__08663__B1 _02029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11668_ net429 net577 _06191_ net300 net1468 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__a32o_1
XFILLER_0_148_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13407_ clknet_leaf_136_clk _00638_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[395\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ net66 _05361_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12211__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12146__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11599_ net428 net579 _06155_ net304 net1533 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08966__A1 final_design.CPU_instr_adr\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07313__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13338_ clknet_leaf_151_clk _00569_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[326\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11970__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13269_ clknet_leaf_28_clk _00500_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[257\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09915__A0 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12514__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11722__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ final_design.cpu.reg_window\[469\] final_design.cpu.reg_window\[501\] net884
+ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07761_ _02708_ _02709_ _02710_ _02711_ net693 net712 vssd1 vssd1 vccd1 vccd1 _02712_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12278__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ _04124_ _04418_ _04417_ net265 vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__o211a_1
X_06712_ final_design.cpu.reg_window\[88\] final_design.cpu.reg_window\[120\] net950
+ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__mux2_1
X_07692_ _01599_ _02513_ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09431_ _03585_ _03589_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__or2_1
X_06643_ _01590_ _01591_ _01592_ _01593_ net788 net794 vssd1 vssd1 vccd1 vccd1 _01594_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11733__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06901__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08329__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09362_ _04158_ _04164_ _02738_ _04133_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_47_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06574_ final_design.cpu.reg_window\[989\] final_design.cpu.reg_window\[1021\] net959
+ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06546__C net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08313_ final_design.cpu.reg_window\[328\] final_design.cpu.reg_window\[360\] net839
+ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07001__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09293_ _02641_ _04088_ _04206_ _04209_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__o211a_1
XANTENNA_11 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08244_ net605 _03192_ _03168_ net541 vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12202__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08175_ final_design.cpu.reg_window\[527\] final_design.cpu.reg_window\[559\] net824
+ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__mux2_1
XANTENNA__12056__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1145_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07126_ _02073_ _02074_ _02075_ _02076_ net783 net802 vssd1 vssd1 vccd1 vccd1 _02077_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_132_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10764__A1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11961__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11895__S net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07057_ net759 _02007_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__nor2_1
XANTENNA__09873__B _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__12505__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07068__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10812__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11196__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ _02906_ _02907_ _02908_ _02909_ net686 net706 vssd1 vssd1 vccd1 vccd1 _02910_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ net85 net1059 vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07613__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09629_ _02868_ _02898_ _04331_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__and3b_1
XANTENNA__11643__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ _06307_ net1459 net992 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12571_ net2127 _06290_ _06286_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__mux2_1
XANTENNA__12441__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_156_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11522_ net2318 net199 net524 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__mux2_1
XANTENNA__07543__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08671__C _01628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ net1306 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_163_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11453_ net239 net2516 net309 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__mux2_1
X_10404_ _03450_ _05181_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__nor2_1
X_14172_ clknet_leaf_81_clk _01346_ net1247 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11384_ net746 _03821_ _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__a21o_1
XANTENNA__10755__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10755__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13123_ clknet_leaf_7_clk _00354_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_10335_ net1490 net1022 net999 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1
+ vccd1 _00092_ sky130_fd_sc_hd__a22o_1
X_13054_ clknet_leaf_19_clk _00285_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_10266_ final_design.uart.BAUD_counter\[24\] _05128_ net809 vssd1 vssd1 vccd1 vccd1
+ _05130_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11704__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ _06207_ net281 net400 net1762 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10197_ final_design.uart.BAUD_counter\[5\] final_design.uart.BAUD_counter\[4\] final_design.uart.BAUD_counter\[8\]
+ final_design.uart.BAUD_counter\[9\] vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__or4b_1
XFILLER_0_17_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09125__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11393__X _06078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13956_ clknet_leaf_107_clk _01187_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[944\]
+ sky130_fd_sc_hd__dfrtp_1
X_12907_ clknet_leaf_133_clk _00145_ net1166 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07231__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13887_ clknet_leaf_137_clk _01118_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[875\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11045__S net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12838_ clknet_leaf_77_clk _00076_ net1254 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07439__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11235__A2 _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12769_ net2566 net808 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_41_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08862__B net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput42 mem_adr_start[15] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_4
Xinput53 mem_adr_start[25] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_1
XFILLER_0_24_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput64 mem_adr_start[6] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_1
XFILLER_0_25_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput75 memory_size[16] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold804 final_design.cpu.reg_window\[663\] vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
Xinput86 memory_size[26] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_2
XANTENNA__10746__A1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold815 final_design.cpu.reg_window\[346\] vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold826 final_design.cpu.reg_window\[507\] vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput97 memory_size[7] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_4
Xhold837 final_design.cpu.reg_window\[505\] vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11943__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold848 final_design.cpu.reg_window\[75\] vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09980_ _03356_ _04706_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_90_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10913__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold859 final_design.cpu.reg_window\[958\] vssd1 vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13286__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08931_ _03758_ _03861_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08862_ net1030 net260 vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__or2_1
XANTENNA__11171__A1 _04825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07813_ _01660_ net621 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__nor2_1
X_08793_ _03680_ _03681_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout186_A _06052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07744_ final_design.cpu.reg_window\[538\] final_design.cpu.reg_window\[570\] net870
+ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06838__A _01785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08529__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07433__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ final_design.cpu.reg_window\[990\] final_design.cpu.reg_window\[1022\] net849
+ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__mux2_1
XANTENNA__12671__B2 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout353_A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ _04331_ _04332_ net449 vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_45_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1095_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__S1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06626_ final_design.cpu.reg_window\[91\] final_design.cpu.reg_window\[123\] net960
+ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09345_ _04057_ _04076_ net473 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06557_ _01453_ _01507_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout520_A net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout618_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_X net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_33_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09276_ net88 _04194_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08264__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06488_ net760 _01430_ net755 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08227_ _03174_ _03175_ _03176_ _03177_ net691 net711 vssd1 vssd1 vccd1 vccd1 _03178_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07850__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1050_X net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08158_ final_design.cpu.reg_window\[399\] final_design.cpu.reg_window\[431\] net826
+ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__mux2_1
XANTENNA__12581__Y _06296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11934__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07109_ final_design.data_from_mem\[12\] net1051 net1008 net1005 vssd1 vssd1 vccd1
+ vccd1 _02060_ sky130_fd_sc_hd__or4_2
X_08089_ _02902_ _03033_ _03037_ _03039_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__a211oi_4
X_10120_ _01370_ _05027_ _05029_ _04999_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[6\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07608__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_42_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10051_ _04654_ _04656_ _04700_ _04748_ _04749_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07461__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12771__2 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__inv_2
X_13810_ clknet_leaf_40_clk _01041_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[798\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13741_ clknet_leaf_139_clk _00972_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[729\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11373__B net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ _05680_ _05676_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__and2b_1
XANTENNA__07213__S0 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13672_ clknet_leaf_117_clk _00903_ net1193 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[660\]
+ sky130_fd_sc_hd__dfrtp_1
X_10884_ _05613_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ final_design.VGA_data_control.state\[0\] final_design.VGA_data_control.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__xor2_2
XFILLER_0_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12554_ _06217_ net346 net323 net2025 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__a22o_1
XANTENNA__09291__A0 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08174__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13797__RESET_B net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11505_ net1740 net227 net526 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12485_ _06145_ net355 net333 net2416 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14224_ final_design.pixel_data vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11436_ net1756 net186 net313 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__mux2_1
XANTENNA__11925__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14155_ clknet_leaf_78_clk _01329_ net1250 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11367_ net748 _03837_ _06054_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ clknet_leaf_44_clk _00337_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_60_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10318_ net1508 net1022 net999 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1
+ vccd1 _00075_ sky130_fd_sc_hd__a22o_1
X_14086_ clknet_leaf_96_clk _01283_ net1229 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11548__B net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11298_ net651 _05994_ _05993_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__a21o_1
XANTENNA__10452__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08149__A2 _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13037_ clknet_leaf_140_clk _00268_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10249_ final_design.uart.BAUD_counter\[18\] _05118_ vssd1 vssd1 vccd1 vccd1 _05119_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_119_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12350__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1140 net1145 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__clkbuf_4
Xfanout1151 net1152 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__clkbuf_4
Xfanout1162 net1163 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__clkbuf_2
Xfanout1173 net1189 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__buf_2
Xfanout1184 net1188 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__clkbuf_4
Xfanout1195 net1196 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08349__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13939_ clknet_leaf_35_clk _01170_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[927\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12653__B2 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07460_ final_design.cpu.reg_window\[896\] final_design.cpu.reg_window\[928\] net951
+ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06411_ final_design.CPU_instr_adr\[4\] vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
X_07391_ _02338_ _02339_ _02340_ _02341_ net785 net803 vssd1 vssd1 vccd1 vccd1 _02342_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11503__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_14_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ _02771_ _03594_ _03599_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__a21boi_1
XANTENNA__07489__A _02185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09282__A0 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10967__A1 _05673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09061_ net631 _03983_ _03985_ _03655_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08012_ net617 _02961_ _02937_ _01937_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold601 final_design.cpu.reg_window\[572\] vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold612 final_design.cpu.reg_window\[42\] vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 final_design.cpu.reg_window\[432\] vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 final_design.cpu.reg_window\[785\] vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 final_design.cpu.reg_window\[49\] vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11392__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold656 final_design.cpu.reg_window\[518\] vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 final_design.cpu.reg_window\[887\] vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09963_ _04851_ _04864_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__xor2_1
XANTENNA__11458__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 final_design.cpu.reg_window\[859\] vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 final_design.cpu.reg_window\[533\] vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_135_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08914_ _02468_ _03856_ _03857_ net629 net259 vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1010_A _06295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ _03558_ _03559_ _03638_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1108_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12341__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08845_ final_design.CPU_instr_adr\[22\] final_design.CPU_instr_adr\[21\] _03795_
+ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout470_A _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_X net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ _03696_ _03726_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__nor2_1
XANTENNA__08259__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06571__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_108_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07016__X _01967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07727_ final_design.cpu.reg_window\[410\] final_design.cpu.reg_window\[442\] net873
+ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout735_A _01493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07658_ _02608_ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06609_ final_design.cpu.reg_window\[732\] final_design.cpu.reg_window\[764\] net954
+ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ net889 _02521_ _02527_ _02533_ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__o32a_4
XTAP_TAPCELL_ROW_153_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11413__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09328_ net322 _04052_ _04246_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_153_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09812__A2 _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ net90 net93 net94 vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__and3_1
XANTENNA__08171__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_117_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12270_ net573 _06200_ net509 net368 net1925 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11907__A0 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout892_X net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ _04744_ net661 vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11383__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07338__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09119__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _02358_ _05838_ net679 vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07682__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10103_ final_design.VGA_data_control.v_count\[0\] _05017_ _05018_ vssd1 vssd1 vccd1
+ vccd1 final_design.vga.v_next_count\[0\] sky130_fd_sc_hd__o21a_1
X_11083_ net91 _05780_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12332__B1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08536__C1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _04950_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__nor2_1
XANTENNA__11686__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08677__B _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11985_ _06187_ net292 net407 net1788 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__a22o_1
XANTENNA__12635__B2 final_design.data_from_mem\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09500__A1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10936_ _05643_ _05647_ _05664_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__or3_1
X_13724_ clknet_leaf_152_clk _00955_ net1117 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[712\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13978__RESET_B net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07801__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10867_ net676 _05584_ _05598_ net977 _05597_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__o221a_1
XANTENNA__10287__X _05143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13655_ clknet_leaf_137_clk _00886_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[643\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10728__A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12399__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12606_ net1437 net1010 net996 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1
+ vccd1 _01299_ sky130_fd_sc_hd__a22o_1
X_13586_ clknet_leaf_42_clk _00817_ net1150 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[574\]
+ sky130_fd_sc_hd__dfrtp_1
X_10798_ _05512_ _05514_ _05531_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12537_ _06200_ net344 net323 net1964 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__a22o_1
XANTENNA__11610__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12468_ _06128_ net353 net333 net2336 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09567__A1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14207_ net1276 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
X_11419_ net2071 net217 net312 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__mux2_1
XANTENNA__12154__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12399_ _06097_ net355 net341 net2290 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__a22o_1
XANTENNA__11374__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14138_ clknet_leaf_76_clk final_design.vga.h_next_count\[7\] net1252 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.VGA_request_address\[1\] sky130_fd_sc_hd__dfrtp_1
X_14069_ clknet_leaf_52_clk _00039_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.uart.receiving
+ sky130_fd_sc_hd__dfrtp_1
X_06960_ _01908_ _01910_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__and2_1
XANTENNA__11126__A1 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06891_ _01838_ _01839_ _01840_ _01841_ net775 net796 vssd1 vssd1 vccd1 vccd1 _01842_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_33_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08630_ _03102_ _03580_ _03579_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__a21o_1
XANTENNA__07976__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08561_ net726 _03511_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__or2_1
X_07512_ _01825_ _02460_ _01790_ _01824_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_18_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07728__S1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08492_ _03439_ _03440_ _03441_ _03442_ net692 net714 vssd1 vssd1 vccd1 vccd1 _03443_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_147_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07443_ _02391_ _02393_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__nand2_2
XFILLER_0_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10638__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07374_ net899 _02318_ _02324_ _02311_ _02312_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_134_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09113_ _02419_ _02424_ net629 vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11601__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout316_A _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09044_ _03973_ _03968_ net258 vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__mux2_1
XANTENNA__07947__A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06851__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09558__A1 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold420 final_design.cpu.reg_window\[981\] vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 final_design.cpu.reg_window\[254\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08114__Y _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11365__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold442 final_design.cpu.reg_window\[766\] vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1225_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold453 final_design.cpu.reg_window\[773\] vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold464 final_design.cpu.reg_window\[680\] vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold475 final_design.cpu.reg_window\[901\] vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold486 final_design.cpu.reg_window\[133\] vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout900 _01437_ vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__buf_4
XANTENNA_fanout685_A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout911 net912 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_4
Xhold497 final_design.cpu.reg_window\[976\] vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout922 net966 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_2
X_09946_ net534 net533 _02325_ net532 net455 net464 vssd1 vssd1 vccd1 vccd1 _04865_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_74_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1013_X net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout933 net966 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_4
Xfanout944 net945 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_4
Xfanout955 net956 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_4
Xfanout966 _01420_ vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__buf_6
Xfanout977 net979 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ net533 net459 _04063_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__a21o_1
Xhold1120 final_design.cpu.reg_window\[816\] vssd1 vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout852_A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout988 _06299_ vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__clkbuf_2
Xfanout999 net1000 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__buf_2
Xhold1131 final_design.cpu.reg_window\[626\] vssd1 vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08533__A2 _03481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10876__B1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 final_design.cpu.reg_window\[631\] vssd1 vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ _03657_ _03778_ _03656_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__a21o_1
Xhold1153 final_design.cpu.reg_window\[312\] vssd1 vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 final_design.cpu.reg_window\[306\] vssd1 vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 final_design.cpu.reg_window\[226\] vssd1 vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1186 final_design.uart.bits_received\[3\] vssd1 vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1197 final_design.uart.BAUD_counter\[7\] vssd1 vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12617__A1 final_design.reqhand.data_from_UART\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08759_ final_design.CPU_instr_adr\[3\] _02330_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _05848_ net595 vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_120_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06585__X _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12747__B net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10721_ _05436_ _05457_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__and2_1
XANTENNA__11651__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13440_ clknet_leaf_35_clk _00671_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[428\]
+ sky130_fd_sc_hd__dfrtp_1
X_10652_ _05389_ _05393_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_125_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13371_ clknet_leaf_136_clk _00602_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[359\]
+ sky130_fd_sc_hd__dfrtp_1
X_10583_ net1488 net1046 net1016 _05328_ vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12322_ net2101 net189 net366 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input79_A memory_size[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09549__A1 _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ net566 _06182_ net505 net372 net1471 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__a32o_1
XFILLER_0_160_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11204_ net432 net583 _05911_ net317 net2121 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__a32o_1
XANTENNA__12553__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11014__C_N net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12184_ net1723 net197 net382 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12953__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ _02358_ net815 net817 vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__or3b_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11066_ net971 _05785_ _05788_ _04042_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06700__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__X _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14106__RESET_B net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ _03627_ _03649_ _03611_ _03617_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__or4bb_1
XANTENNA__10331__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06630__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12608__B2 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12084__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11968_ _06170_ net287 net405 net1526 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13707_ clknet_leaf_16_clk _00938_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[695\]
+ sky130_fd_sc_hd__dfrtp_1
X_10919_ _05647_ _05648_ net2554 net1043 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12149__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11899_ net208 net2137 net275 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__mux2_1
XANTENNA__10458__A _02570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13638_ clknet_leaf_170_clk _00869_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[626\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13569_ clknet_leaf_157_clk _00800_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[557\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11595__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07767__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07090_ final_design.cpu.reg_window\[204\] final_design.cpu.reg_window\[236\] net927
+ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12544__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09800_ _03563_ _04718_ _03391_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09960__A1 _04871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout207 net208 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__buf_2
Xfanout218 _05928_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10921__A net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout229 _05864_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_2
X_07992_ final_design.cpu.reg_window\[80\] final_design.cpu.reg_window\[112\] net879
+ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06943_ _01890_ _01891_ _01892_ _01893_ net775 net796 vssd1 vssd1 vccd1 vccd1 _01894_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06610__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09731_ _04220_ _04408_ _04648_ _04649_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09662_ net486 _04578_ _04579_ _04580_ _04294_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__a32o_1
X_06874_ _01815_ _01823_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_2_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08613_ _03391_ _03563_ _03562_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__a21o_1
X_09593_ _02770_ _04281_ _04168_ _02705_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_141_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout266_A net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13829__RESET_B net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08544_ final_design.cpu.reg_window\[1\] final_design.cpu.reg_window\[33\] net850
+ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07441__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11471__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11283__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08475_ _03359_ _03425_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout433_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1175_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07426_ final_design.cpu.reg_window\[833\] final_design.cpu.reg_window\[865\] net936
+ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13411__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11898__S net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08126__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07357_ final_design.cpu.reg_window\[195\] final_design.cpu.reg_window\[227\] net945
+ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__mux2_1
XANTENNA__10389__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08272__S net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07288_ net895 _02238_ _02227_ _02221_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ final_design.CPU_instr_adr\[12\] net1026 _03956_ _03958_ vssd1 vssd1 vccd1
+ vccd1 _00223_ sky130_fd_sc_hd__a22o_1
XANTENNA__11199__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12535__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold250 final_design.cpu.reg_window\[453\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07637__S0 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09400__B1 _04301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold261 final_design.cpu.reg_window\[95\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 final_design.cpu.reg_window\[457\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold283 final_design.cpu.reg_window\[140\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__A1 _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold294 final_design.cpu.reg_window\[169\] vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout730 net732 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_6
Xfanout741 net742 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07616__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09929_ _04178_ _04829_ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__or3b_1
Xfanout752 net753 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout763 net764 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout774 net776 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__buf_4
Xfanout785 net787 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08506__A2 _03450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout796 net798 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_4
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12940_ clknet_leaf_67_clk _00178_ net1223 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_161_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07562__D net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11510__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10977__S net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ clknet_leaf_79_clk _00109_ net1251 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11822_ net214 net2266 net266 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08447__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07351__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11381__B net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11274__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ net204 net2275 net416 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10704_ net1015 _05442_ _05443_ net1041 net1385 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__a32o_1
XFILLER_0_154_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09482__A3 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11684_ net574 net421 _06200_ net295 net1690 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__a32o_1
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ final_design.CPU_instr_adr\[9\] _05377_ net1069 vssd1 vssd1 vccd1 vccd1 _05378_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13423_ clknet_leaf_97_clk _00654_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[411\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_141_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08690__B net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload109 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__clkinvlp_4
X_13354_ clknet_leaf_3_clk _00585_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[342\]
+ sky130_fd_sc_hd__dfrtp_1
X_10566_ net96 final_design.VGA_adr\[4\] vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12305_ net1812 net220 net365 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__mux2_1
X_13285_ clknet_leaf_18_clk _00516_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[273\]
+ sky130_fd_sc_hd__dfrtp_1
X_10497_ _05233_ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__or2_1
XANTENNA__12526__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12236_ net573 _06166_ net509 net373 net1503 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__a32o_1
X_14199__1268 vssd1 vssd1 vccd1 vccd1 _14199__1268/HI net1268 sky130_fd_sc_hd__conb_1
XANTENNA__10001__A1 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12167_ net2146 net226 net382 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__mux2_1
XANTENNA__12432__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11118_ final_design.uart.bits_received\[0\] final_design.uart.bits_received\[1\]
+ final_design.uart.bits_received\[2\] final_design.uart.bits_received\[3\] vssd1
+ vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__a31o_1
XANTENNA__11556__B net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09307__A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12098_ net1914 net226 net390 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__mux2_1
XANTENNA__10460__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ _01387_ _05772_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__nor2_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
X_06590_ _01536_ _01539_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__nand2_1
XANTENNA__10068__A1 _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09042__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08356__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11804__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08260_ _03207_ _03208_ _03209_ _03210_ net690 net710 vssd1 vssd1 vccd1 vccd1 _03211_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_942 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07211_ final_design.cpu.reg_window\[456\] final_design.cpu.reg_window\[488\] net920
+ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08191_ final_design.cpu.reg_window\[78\] final_design.cpu.reg_window\[110\] net844
+ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11511__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07142_ _01468_ net747 net887 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08092__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__B2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06605__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08984__A2 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07073_ _02020_ _02021_ _02022_ _02023_ net777 net797 vssd1 vssd1 vccd1 vccd1 _02024_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12517__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08292__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ final_design.cpu.reg_window\[529\] final_design.cpu.reg_window\[561\] net827
+ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__mux2_1
XANTENNA__08121__A _02030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09714_ net72 _04184_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__nand2_1
X_06926_ final_design.cpu.reg_window\[530\] final_design.cpu.reg_window\[562\] net901
+ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__mux2_1
XANTENNA__07960__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06857_ net762 _01807_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__nor2_1
X_09645_ _04218_ _04563_ _04556_ net264 _04558_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_97_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout550_A _01880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08775__B _02186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09576_ _03295_ _03569_ _03576_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06788_ final_design.cpu.reg_window\[534\] final_design.cpu.reg_window\[566\] net902
+ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__mux2_1
XANTENNA__08267__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11256__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08527_ final_design.cpu.reg_window\[514\] final_design.cpu.reg_window\[546\] net865
+ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1080_X net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08458_ final_design.cpu.reg_window\[708\] final_design.cpu.reg_window\[740\] net858
+ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11008__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07409_ _01484_ _02358_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_137_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08389_ net718 _03333_ net730 vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11559__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11421__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10420_ net1574 net1047 _05193_ net248 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10351_ net2 net1037 net1020 final_design.data_from_mem\[0\] vssd1 vssd1 vccd1 vccd1
+ _00104_ sky130_fd_sc_hd__o22a_1
XFILLER_0_143_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12508__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06986__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13070_ clknet_leaf_116_clk _00301_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_10282_ net2496 _05138_ net810 vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout972_X net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12021_ _06223_ net293 net403 net2122 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10561__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_163_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08669__C _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09127__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout571 net572 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_4
Xfanout582 _05868_ vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_4
X_13972_ clknet_leaf_101_clk _01203_ net1188 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[960\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout593 net594 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11495__A0 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ clknet_leaf_110_clk _00161_ net1214 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12854_ clknet_leaf_82_clk _00092_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08177__S net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13333__RESET_B net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11247__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11805_ net2355 net415 net292 _06061_ vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08663__A1 _01999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11736_ net230 net2474 net418 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10736__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11667_ net176 net639 vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13406_ clknet_leaf_22_clk _00637_ net1127 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[394\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10618_ net66 _05361_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11598_ net178 net643 vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__and2_2
XFILLER_0_148_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08966__A2 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10549_ final_design.CPU_instr_adr\[5\] _05277_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13337_ clknet_leaf_164_clk _00568_ net1085 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[325\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13268_ clknet_leaf_103_clk _00499_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[256\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09915__A1 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12219_ net567 _06147_ net505 net376 net2400 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__a32o_1
X_13199_ clknet_leaf_94_clk _00430_ net1226 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[187\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07256__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11722__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07760_ final_design.cpu.reg_window\[408\] final_design.cpu.reg_window\[440\] net868
+ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__mux2_1
XANTENNA__08026__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06711_ _01658_ _01660_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07691_ _02543_ _02544_ _02637_ _02639_ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11506__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09430_ net499 _04348_ _04231_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__o21bai_1
X_06642_ final_design.cpu.reg_window\[539\] final_design.cpu.reg_window\[571\] net960
+ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__mux2_1
XANTENNA__06901__A1 _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13074__RESET_B net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08329__S1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ _04046_ _04255_ _04256_ _04279_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_47_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06573_ final_design.cpu.reg_window\[797\] final_design.cpu.reg_window\[829\] net959
+ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13003__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10349__C net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08312_ _02186_ net605 vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11789__B2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06546__D _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09292_ net559 net558 net556 net555 net460 net470 vssd1 vssd1 vccd1 vccd1 _04211_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07001__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _01558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08243_ net605 _03192_ _03168_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10461__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__A _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12738__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A _05864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08174_ final_design.cpu.reg_window\[591\] final_design.cpu.reg_window\[623\] net824
+ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07125_ final_design.cpu.reg_window\[139\] final_design.cpu.reg_window\[171\] net937
+ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10933__X _05662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1040_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1138_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07056_ _02003_ _02004_ _02005_ _02006_ net777 net797 vssd1 vssd1 vccd1 vccd1 _02007_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08550__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09873__C _04308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XANTENNA__09906__A1 _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07068__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07166__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11196__B net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ final_design.cpu.reg_window\[401\] final_design.cpu.reg_window\[433\] net836
+ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09234__X _04153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06909_ final_design.cpu.reg_window\[402\] final_design.cpu.reg_window\[434\] net902
+ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout932_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ final_design.cpu.reg_window\[343\] final_design.cpu.reg_window\[375\] net852
+ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__mux2_1
XANTENNA__11416__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09628_ _02898_ _04331_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11229__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ _04452_ _04455_ _04477_ _04425_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_clk_X clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14198__1267 vssd1 vssd1 vccd1 vccd1 _14198__1267/HI net1267 sky130_fd_sc_hd__conb_1
X_12570_ final_design.uart.receiving final_design.uart.working_data\[5\] vssd1 vssd1
+ vccd1 vccd1 _06290_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ net1918 net201 net524 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06751__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14240_ net1305 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XANTENNA__08671__D _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11452_ net239 net647 vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10403_ net1733 net1048 _05184_ net250 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14171_ clknet_leaf_81_clk _01345_ net1255 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09070__A1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11383_ net668 _03815_ net741 vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input61_A mem_adr_start[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ net1525 net1024 net1001 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1
+ vccd1 _00091_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ clknet_leaf_30_clk _00353_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08460__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13053_ clknet_leaf_12_clk _00284_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10265_ final_design.uart.BAUD_counter\[24\] _05128_ vssd1 vssd1 vccd1 vccd1 _05129_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09128__Y _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11704__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ _06206_ net285 net401 net2006 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10196_ final_design.uart.BAUD_counter\[11\] final_design.uart.BAUD_counter\[10\]
+ final_design.uart.bits_received\[2\] final_design.uart.bits_received\[3\] vssd1
+ vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08008__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout390 net391 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09125__A2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13955_ clknet_leaf_6_clk _01186_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[943\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12906_ clknet_leaf_133_clk _00144_ net1166 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07231__S1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886_ clknet_leaf_146_clk _01117_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[874\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12837_ clknet_leaf_77_clk _00075_ net1253 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12768_ final_design.VGA_adr\[8\] net808 _06402_ net967 vssd1 vssd1 vccd1 vccd1 _01355_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06944__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10757__A2_N net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11719_ net190 net636 vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__and2_1
XANTENNA__11640__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12157__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10443__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12699_ final_design.VGA_data_control.v_count\[5\] _06339_ vssd1 vssd1 vccd1 vccd1
+ _06340_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 mem_adr_start[16] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_2
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput54 mem_adr_start[26] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08939__A2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput65 mem_adr_start[7] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09061__A1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold805 final_design.cpu.reg_window\[397\] vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
Xinput76 memory_size[17] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_2
Xhold816 final_design.VGA_data_control.data_to_VGA\[28\] vssd1 vssd1 vccd1 vccd1 net2169
+ sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 memory_size[27] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput98 memory_size[8] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_4
Xhold827 final_design.cpu.reg_window\[333\] vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 final_design.cpu.reg_window\[662\] vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 final_design.cpu.reg_window\[83\] vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10913__B _05642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ _01789_ _02463_ _01759_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12499__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ _03802_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07375__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07812_ _02750_ _02751_ _02762_ net892 vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a22oi_4
X_08792_ _03688_ _03732_ _03742_ _03687_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__and4b_1
XFILLER_0_74_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07743_ final_design.cpu.reg_window\[602\] final_design.cpu.reg_window\[634\] net870
+ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12120__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09667__A3 _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_A _06081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ final_design.cpu.reg_window\[798\] final_design.cpu.reg_window\[830\] net850
+ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__mux2_1
X_09413_ _02804_ _04330_ _04131_ _02900_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__o211ai_1
X_06625_ _01572_ _01573_ _01574_ _01575_ net788 net806 vssd1 vssd1 vccd1 vccd1 _01576_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout346_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06556_ net749 _01497_ net672 _01506_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__a211o_2
X_09344_ _04261_ _04262_ net498 _04097_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__a211o_1
XANTENNA__12423__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09275_ net86 net87 _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__or3_1
XFILLER_0_157_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06487_ net899 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout513_A _06259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1255_A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06733__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08226_ final_design.cpu.reg_window\[139\] final_design.cpu.reg_window\[171\] net856
+ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14043__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07850__A2 _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08157_ final_design.cpu.reg_window\[463\] final_design.cpu.reg_window\[495\] net826
+ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_X net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07108_ net896 _02051_ _02057_ _02044_ _02045_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__a32o_2
XFILLER_0_28_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07063__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08088_ _01718_ _02839_ _02864_ _02868_ _03038_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout882_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07039_ final_design.cpu.reg_window\[526\] final_design.cpu.reg_window\[558\] net935
+ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__mux2_1
XANTENNA__11000__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ _04919_ _04921_ _04922_ _04968_ _04476_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__o2111a_1
XANTENNA__08012__C1 _01937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__A2 _05143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07461__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13740_ clknet_leaf_125_clk _00971_ net1196 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[728\]
+ sky130_fd_sc_hd__dfrtp_1
X_10952_ net84 _05651_ _05679_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__a21o_1
XANTENNA__07213__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10673__A1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13671_ clknet_leaf_9_clk _00902_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[659\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11870__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ _05590_ _05593_ _05611_ _05612_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_123_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12622_ final_design.VGA_data_control.state\[1\] _01402_ final_design.VGA_data_control.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08455__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12414__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09815__B1 _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ _06216_ net343 net323 net2395 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__a22o_1
XANTENNA__11622__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09291__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11504_ net2487 net241 net526 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12484_ _06144_ net345 net331 net2077 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14223_ final_design.v_out vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11669__X _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11435_ net1943 net188 net313 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14154_ clknet_leaf_78_clk _01328_ net1255 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11366_ net668 _03832_ net740 vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__o21a_1
XANTENNA__11388__Y _06074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06703__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10317_ net1524 net1023 net999 final_design.data_from_mem\[2\] vssd1 vssd1 vccd1
+ vccd1 _00074_ sky130_fd_sc_hd__a22o_1
X_13105_ clknet_leaf_109_clk _00336_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[93\]
+ sky130_fd_sc_hd__dfrtp_1
X_14085_ clknet_leaf_71_clk _01282_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11297_ final_design.data_from_mem\[18\] net235 net233 vssd1 vssd1 vccd1 vccd1 _05994_
+ sky130_fd_sc_hd__a21o_2
X_10248_ _05118_ net809 _05117_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__and3b_1
X_13036_ clknet_leaf_123_clk _00267_ net1191 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1130 net1132 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__clkbuf_4
Xfanout1141 net1145 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__clkbuf_2
X_10179_ final_design.uart.BAUD_counter\[25\] final_design.uart.BAUD_counter\[24\]
+ final_design.uart.BAUD_counter\[27\] final_design.uart.BAUD_counter\[26\] vssd1
+ vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__or4_1
Xfanout1152 net1153 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12440__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1163 net1164 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1174 net1177 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__clkbuf_4
Xfanout1185 net1188 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__buf_2
XANTENNA__07534__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11564__B net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1196 net1217 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13938_ clknet_leaf_41_clk _01169_ net1150 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[926\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_8__f_clk_X clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11861__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13869_ clknet_leaf_127_clk _01100_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[857\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06410_ final_design.CPU_instr_adr\[12\] vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11580__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07390_ final_design.cpu.reg_window\[130\] final_design.cpu.reg_window\[162\] net939
+ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08365__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12405__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06674__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07489__B _02186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10416__B2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09282__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09060_ _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09985__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08011_ _01939_ net609 vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10924__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold602 final_design.cpu.reg_window\[365\] vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold613 final_design.cpu.reg_window\[426\] vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 final_design.cpu.reg_window\[999\] vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold635 final_design.cpu.reg_window\[270\] vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold646 final_design.cpu.reg_window\[893\] vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 final_design.cpu.reg_window\[225\] vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold668 final_design.cpu.reg_window\[132\] vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ net90 _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_38_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold679 final_design.cpu.reg_window\[81\] vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08913_ _03768_ _03770_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__xnor2_1
X_14197__1266 vssd1 vssd1 vccd1 vccd1 _14197__1266/HI net1266 sky130_fd_sc_hd__conb_1
X_09893_ _03558_ _03559_ _03638_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout296_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__C1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ final_design.CPU_instr_adr\[20\] _03794_ vssd1 vssd1 vccd1 vccd1 _03795_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_85_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10352__B1 _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08775_ final_design.CPU_instr_adr\[8\] _02186_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout463_A _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07726_ final_design.cpu.reg_window\[474\] final_design.cpu.reg_window\[506\] net873
+ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout251_X net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout630_A _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07657_ _02605_ _02607_ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11490__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout728_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06608_ net763 _01558_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_101_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07588_ net719 _02538_ net889 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_153_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06539_ _01464_ _01475_ _01483_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__nor3_2
XANTENNA__10407__B2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09327_ _02641_ _03607_ _04051_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_153_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08076__A2 _03022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1160_X net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09258_ net733 _04127_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__or3_2
XFILLER_0_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08209_ net889 _03141_ _03147_ _03153_ _03159_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__o32a_2
X_09189_ net485 _04054_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11220_ net652 _05925_ _05924_ _05142_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11649__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11151_ net655 net228 vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__and2_1
XANTENNA__07682__S1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ final_design.VGA_data_control.v_count\[0\] _05017_ _05007_ vssd1 vssd1 vccd1
+ vccd1 _05018_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_105_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11082_ _05780_ _05802_ _05803_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__nor3_1
XANTENNA__13106__RESET_B net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ _04330_ _04951_ net449 vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11665__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09406__Y _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06759__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11984_ _06186_ net291 net406 net1646 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__a22o_1
X_13723_ clknet_leaf_155_clk _00954_ net1115 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[711\]
+ sky130_fd_sc_hd__dfrtp_1
X_10935_ _05662_ net243 vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ clknet_leaf_124_clk _00885_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[642\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08185__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10866_ final_design.CPU_instr_adr\[20\] net1013 _05595_ net1054 vssd1 vssd1 vccd1
+ vccd1 _05598_ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06494__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ net1395 net1009 net995 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1
+ vccd1 _01298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09264__A1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13585_ clknet_leaf_107_clk _00816_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[573\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10797_ _05512_ _05514_ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12536_ _06199_ net343 net323 net2391 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__a22o_1
XANTENNA__07814__A2 _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13947__RESET_B net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12467_ _06127_ net355 net333 net2068 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__a22o_1
XANTENNA__12435__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14206_ net1275 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07529__S net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11418_ net1754 net219 net311 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__mux2_1
XANTENNA__12020__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09567__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12398_ _06096_ net350 net340 net2333 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11374__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14137_ clknet_leaf_75_clk final_design.vga.h_next_count\[6\] net1253 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.VGA_request_address\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11349_ net434 net586 _06039_ net317 net1767 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14068_ clknet_leaf_52_clk _00038_ net1153 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter_state
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11126__A2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12170__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ clknet_leaf_156_clk _00250_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_06890_ final_design.cpu.reg_window\[915\] final_design.cpu.reg_window\[947\] net908
+ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08560_ _03507_ _03508_ _03509_ _03510_ net689 net701 vssd1 vssd1 vccd1 vccd1 _03511_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12087__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07189__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10637__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07511_ _01824_ _02461_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11834__A0 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10637__B2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08491_ final_design.cpu.reg_window\[899\] final_design.cpu.reg_window\[931\] net861
+ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11514__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07442_ _01484_ net815 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_174_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07373_ net771 _02323_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09112_ _03715_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09043_ _02444_ net631 _03969_ _03972_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__a31o_1
XFILLER_0_154_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout211_A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13617__RESET_B net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold410 final_design.cpu.reg_window\[586\] vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12011__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold421 final_design.cpu.reg_window\[87\] vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 final_design.cpu.reg_window\[650\] vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 final_design.cpu.reg_window\[165\] vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11365__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold454 final_design.cpu.reg_window\[729\] vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1120_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 final_design.cpu.reg_window\[906\] vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold476 final_design.cpu.reg_window\[591\] vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold487 final_design.cpu.reg_window\[596\] vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1218_A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout901 net903 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__clkbuf_4
Xhold498 final_design.cpu.reg_window\[975\] vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
X_09945_ net734 _04863_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__nor2_1
Xfanout912 net922 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout923 net924 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12314__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout934 net935 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08518__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net966 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_4
Xfanout956 net966 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__buf_2
Xfanout967 _05039_ vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ net538 net537 net536 net534 net454 net463 vssd1 vssd1 vccd1 vccd1 _04795_
+ sky130_fd_sc_hd__mux4_1
Xfanout978 net979 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_4
Xhold1110 final_design.cpu.reg_window\[117\] vssd1 vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 _06299_ vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__buf_2
Xhold1121 final_design.cpu.reg_window\[256\] vssd1 vssd1 vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 final_design.cpu.reg_window\[622\] vssd1 vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10876__A1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08827_ _01358_ _01538_ _03777_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a21oi_1
Xhold1143 final_design.uart.BAUD_counter\[30\] vssd1 vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 final_design.cpu.reg_window\[638\] vssd1 vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1165 final_design.cpu.reg_window\[821\] vssd1 vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1176 final_design.reqhand.instruction\[6\] vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 net124 vssd1 vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12078__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08758_ final_design.CPU_instr_adr\[3\] _02330_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__and2_1
Xhold1198 final_design.uart.BAUD_counter\[4\] vssd1 vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07902__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11825__A0 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07709_ _02656_ _02657_ _02658_ _02659_ net696 net715 vssd1 vssd1 vccd1 vccd1 _02660_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08689_ net622 _03549_ _03523_ _02419_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__a211o_1
XFILLER_0_166_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06927__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11424__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12093__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _05438_ _05441_ _05457_ _05436_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07203__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _05391_ _05392_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09246__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10582_ _05309_ _05326_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__xnor2_1
X_13370_ clknet_leaf_163_clk _00601_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[358\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12250__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09797__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12321_ net2104 net191 net366 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12252_ net596 _06181_ net519 net375 net1923 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__a32o_1
XANTENNA__12002__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11203_ net656 net244 vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__and2_1
XANTENNA__09954__C1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12183_ net1891 net199 net380 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ net815 net817 _02359_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__and3b_4
X_11065_ _01358_ _03821_ net1072 vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__mux2_1
XANTENNA__07084__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ net264 _04928_ _04934_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10867__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12993__RESET_B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10867__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12069__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14146__RESET_B net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09485__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ _06169_ net284 net405 net1625 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ clknet_leaf_2_clk _00937_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[694\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10918_ _05624_ _05645_ _05646_ net1018 vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11898_ net210 net2158 net275 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10458__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_134_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13637_ clknet_leaf_4_clk _00868_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[625\]
+ sky130_fd_sc_hd__dfrtp_1
X_10849_ _05559_ _05564_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__or3_1
X_14196__1265 vssd1 vssd1 vccd1 vccd1 _14196__1265/HI net1265 sky130_fd_sc_hd__conb_1
XFILLER_0_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12796__27 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__inv_2
XFILLER_0_66_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07248__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11044__B2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12241__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13568_ clknet_leaf_37_clk _00799_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[556\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08996__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11595__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12519_ _06181_ net359 net330 net1773 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__a22o_1
XANTENNA__10474__A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12165__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13499_ clknet_leaf_153_clk _00730_ net1116 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[487\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_149_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06471__A1 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07259__S net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout208 _05965_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
Xfanout219 _05921_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_2
XFILLER_0_10_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07991_ _02938_ _02939_ _02940_ _02941_ net696 net715 vssd1 vssd1 vccd1 vccd1 _02942_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10921__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11509__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09730_ net497 _04113_ _04268_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__or3_1
X_06942_ final_design.cpu.reg_window\[145\] final_design.cpu.reg_window\[177\] net910
+ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09661_ net486 _04225_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__nor2_1
X_06873_ _01815_ _01823_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_2_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08612_ _02294_ net499 vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__nor2_1
X_09592_ net736 _04502_ _04508_ _04482_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_141_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09503__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08543_ final_design.cpu.reg_window\[65\] final_design.cpu.reg_window\[97\] net850
+ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__mux2_1
XANTENNA__11807__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09476__A1 _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__A3 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout259_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11283__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12480__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ _03387_ _03389_ _03420_ _03422_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__o22a_1
XFILLER_0_148_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07425_ net760 _02369_ net755 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout426_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1168_A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08553__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ final_design.cpu.reg_window\[3\] final_design.cpu.reg_window\[35\] net942
+ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__mux2_1
XANTENNA__08436__C1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07287_ _02232_ _02237_ net766 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__mux2_1
XANTENNA__10384__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09026_ net257 _03957_ net1027 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout795_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold240 final_design.cpu.reg_window\[588\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold251 final_design.cpu.reg_window\[44\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold262 final_design.cpu.reg_window\[858\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07637__S1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold273 final_design.uart.BAUD_counter\[25\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10010__A2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold284 final_design.cpu.reg_window\[690\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 final_design.cpu.reg_window\[756\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout962_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 net724 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout731 net732 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11419__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout742 _01491_ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__buf_2
X_09928_ _04843_ _04845_ net733 _04831_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a211o_2
Xfanout753 _01476_ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_2
Xfanout764 net765 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_4
Xfanout775 net776 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_4
XFILLER_0_99_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout786 net787 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__buf_4
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout797 net798 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__buf_4
X_09859_ net541 net540 net539 net538 net454 net463 vssd1 vssd1 vccd1 vccd1 _04778_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ clknet_leaf_79_clk _00108_ net1250 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11821_ net215 net1849 net266 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__mux2_1
XANTENNA__12066__A3 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11274__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07204__Y _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12471__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11752_ net221 net2274 net418 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10703_ _05438_ _05441_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__or2_1
X_11683_ net238 net635 vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input91_A memory_size[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13422_ clknet_leaf_114_clk _00653_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[410\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10634_ _05351_ _05376_ _05371_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__o21a_1
XANTENNA__12223__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06772__A _01718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08463__S net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11577__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08978__B1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13353_ clknet_leaf_88_clk _00584_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[341\]
+ sky130_fd_sc_hd__dfrtp_1
X_10565_ net96 final_design.VGA_adr\[4\] vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12304_ net1919 net244 net364 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__mux2_1
XANTENNA__07650__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13284_ clknet_leaf_100_clk _00515_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[272\]
+ sky130_fd_sc_hd__dfrtp_1
X_10496_ _05244_ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__nand2b_1
XANTENNA__11329__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12235_ net568 _06165_ net508 net372 net1578 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__a32o_1
XANTENNA__08699__A _02510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09147__X _04066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__Y _06081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12166_ net1941 net241 net382 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ final_design.uart.bits_received\[2\] _05830_ _05831_ _05834_ vssd1 vssd1
+ vccd1 vccd1 _00207_ sky130_fd_sc_hd__a22o_1
X_12097_ net2011 net241 net390 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048_ net677 _05758_ _05771_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__o21ai_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07542__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11572__B net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12999_ net1341 _00230_ net1159 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09610__X _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07210_ final_design.cpu.reg_window\[264\] final_design.cpu.reg_window\[296\] net921
+ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12214__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08190_ net719 _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07141_ _01488_ net738 _01820_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__or3b_1
XFILLER_0_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07072_ final_design.cpu.reg_window\[909\] final_design.cpu.reg_window\[941\] net915
+ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_144_Left_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10932__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09394__B1 _04231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08292__S1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07974_ final_design.cpu.reg_window\[593\] final_design.cpu.reg_window\[625\] net827
+ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09713_ net735 _04631_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__or2_1
XANTENNA__07018__A _01966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06925_ final_design.cpu.reg_window\[594\] final_design.cpu.reg_window\[626\] net901
+ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout376_A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ _04342_ _04561_ _04562_ _04222_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__o211a_1
X_06856_ _01803_ _01804_ _01805_ _01806_ net787 net803 vssd1 vssd1 vccd1 vccd1 _01807_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06857__A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12578__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07452__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_153_Left_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09575_ net263 _04484_ _04493_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__and3_1
XFILLER_0_139_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06787_ final_design.cpu.reg_window\[598\] final_design.cpu.reg_window\[630\] net902
+ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout543_A _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08526_ final_design.cpu.reg_window\[578\] final_design.cpu.reg_window\[610\] net865
+ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08657__C1 _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout710_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08457_ _03404_ _03405_ _03406_ _03407_ net691 net711 vssd1 vssd1 vccd1 vccd1 _03408_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout331_X net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_X net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13632__RESET_B net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07408_ final_design.data_from_mem\[9\] net981 _02357_ vssd1 vssd1 vccd1 vccd1 _02359_
+ sky130_fd_sc_hd__o21ai_2
XANTENNA__12205__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08283__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ net725 _03338_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11559__A2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07339_ final_design.cpu.reg_window\[580\] final_design.cpu.reg_window\[612\] net939
+ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_162_Left_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10350_ wb_manage.BUSY_O net1039 wb_manage.prev_BUSY_O vssd1 vssd1 vccd1 vccd1 _05171_
+ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_115_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09009_ net257 _03940_ _03941_ _03942_ net1026 vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10281_ final_design.uart.BAUD_counter\[30\] _05138_ vssd1 vssd1 vccd1 vccd1 _05139_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_143_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10842__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_3_0_clk_X clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__A0 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _06222_ net291 net402 net1837 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__a22o_1
XANTENNA__07627__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09408__A _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout965_X net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08312__A _02186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09127__B _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 _01880_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_2
X_14195__1264 vssd1 vssd1 vccd1 vccd1 _14195__1264/HI net1264 sky130_fd_sc_hd__conb_1
Xfanout572 net576 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_2
Xfanout583 net585 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_2
X_13971_ clknet_leaf_35_clk _01202_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[959\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout594 net597 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_171_Left_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12922_ clknet_leaf_11_clk _00160_ net1092 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12692__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08896__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08458__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07362__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12853_ clknet_leaf_86_clk _00091_ net1235 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11247__A1 _04639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11804_ net2287 net414 net291 _06053_ vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__a22o_1
XANTENNA__08405__A_N net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11798__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11735_ net816 _05846_ _05867_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08663__A2 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input94_X net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11666_ net428 net579 _06190_ net300 net1470 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12774__5_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13405_ clknet_leaf_31_clk _00636_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[393\]
+ sky130_fd_sc_hd__dfrtp_1
X_10617_ net676 _05348_ _05360_ net979 _05359_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__o221a_1
XFILLER_0_148_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11597_ net437 net592 _06154_ net306 net1990 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__a32o_1
XANTENNA__12211__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13336_ clknet_leaf_138_clk _00567_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[324\]
+ sky130_fd_sc_hd__dfrtp_1
X_10548_ _05293_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__or2_1
Xclkbuf_4_5__f_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__11970__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12443__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13267_ clknet_leaf_32_clk _00498_ net1129 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[255\]
+ sky130_fd_sc_hd__dfrtp_1
X_10479_ net47 _05223_ _05225_ _05227_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__nand4_1
XFILLER_0_122_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12218_ net595 _06146_ net519 net379 net1879 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__a32o_1
XANTENNA__09318__A net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ clknet_leaf_115_clk _00429_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[186\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11722__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ net199 net2449 net384 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08026__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__A3 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ _01658_ _01660_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12683__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07690_ _02640_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06641_ final_design.cpu.reg_window\[603\] final_design.cpu.reg_window\[635\] net960
+ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ _04056_ _04278_ _04274_ net264 vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_47_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06572_ final_design.cpu.reg_window\[861\] final_design.cpu.reg_window\[893\] net959
+ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11789__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08311_ _03259_ _03260_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09291_ net559 net558 net460 vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11522__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_13 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08242_ _02097_ net619 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10461__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10646__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08173_ final_design.cpu.reg_window\[655\] final_design.cpu.reg_window\[687\] net824
+ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08406__A2 _03352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12202__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ final_design.cpu.reg_window\[203\] final_design.cpu.reg_window\[235\] net937
+ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__mux2_1
XANTENNA__11410__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07055_ final_design.cpu.reg_window\[397\] final_design.cpu.reg_window\[429\] net914
+ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__mux2_1
XANTENNA__11961__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__clkbuf_4
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__clkbuf_4
X_12780__11 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__inv_2
XFILLER_0_30_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07447__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08132__A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout493_A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1200_A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ final_design.cpu.reg_window\[465\] final_design.cpu.reg_window\[497\] net836
+ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout660_A _05143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout758_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ final_design.cpu.reg_window\[466\] final_design.cpu.reg_window\[498\] net903
+ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__mux2_1
X_07888_ _01722_ net607 vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__nand2_1
XANTENNA__07182__S net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09627_ _04046_ _04545_ _04543_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__a21o_1
X_06839_ _01785_ _01788_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ _04452_ _04455_ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a21boi_1
XANTENNA__12426__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08509_ final_design.cpu.reg_window\[450\] final_design.cpu.reg_window\[482\] net860
+ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ net486 _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11432__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11520_ net1845 net204 net524 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08307__A _02157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06751__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire225 _05897_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
XFILLER_0_136_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ net226 net2489 net309 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10402_ _03481_ _05181_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__nor2_1
X_14170_ clknet_leaf_81_clk _01344_ net1247 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11401__A1 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11382_ net435 net589 _06068_ net317 net1727 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__a32o_1
XFILLER_0_61_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13121_ clknet_leaf_159_clk _00352_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10333_ net1548 net1024 net1001 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1
+ vccd1 _00090_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07357__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input54_A mem_adr_start[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ clknet_leaf_149_clk _00283_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_10264_ _05128_ net809 _05127_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__and3b_1
X_12003_ _06205_ net288 net402 net2116 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__a22o_1
XANTENNA__11704__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10195_ _05082_ _05083_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08008__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13__f_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_6
Xfanout391 _06265_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_4
X_13954_ clknet_leaf_29_clk _01185_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[942\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12665__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08188__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ clknet_leaf_131_clk _00143_ net1166 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13885_ clknet_leaf_14_clk _01116_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[873\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12836_ clknet_leaf_75_clk _00074_ net1253 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12417__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ _01369_ _01398_ _06383_ _06398_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12438__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08636__A2 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06647__A1 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11640__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11718_ net429 net578 _06217_ net296 net2172 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__a32o_1
XANTENNA__10443__A2 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12698_ _01368_ _06334_ _06336_ _06337_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__o31a_2
XANTENNA__08217__A _02097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_11649_ net194 net638 vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_1
XFILLER_0_71_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput44 mem_adr_start[17] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput55 mem_adr_start[27] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput66 mem_adr_start[8] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06960__A _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput77 memory_size[18] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_2
Xhold806 final_design.cpu.reg_window\[1008\] vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 final_design.cpu.reg_window\[1003\] vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 memory_size[28] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10746__A3 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold828 final_design.cpu.reg_window\[135\] vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11578__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13319_ clknet_leaf_16_clk _00550_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[307\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11943__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput99 memory_size[9] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_2
XFILLER_0_161_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12173__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold839 final_design.cpu.reg_window\[347\] vssd1 vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07267__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09048__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11156__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08860_ final_design.CPU_instr_adr\[30\] _03801_ vssd1 vssd1 vccd1 vccd1 _03810_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09990__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ _02756_ _02761_ net721 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__mux2_1
X_08791_ _03683_ _03685_ _03686_ _03739_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__and4_1
XFILLER_0_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11517__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07742_ final_design.cpu.reg_window\[666\] final_design.cpu.reg_window\[698\] net870
+ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08098__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08324__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10131__A1 final_design.VGA_data_control.v_count\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07673_ final_design.cpu.reg_window\[862\] final_design.cpu.reg_window\[894\] net849
+ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__mux2_1
X_09412_ _02802_ _02834_ _04330_ _02900_ _02800_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__a311o_1
XANTENNA__12408__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06624_ final_design.cpu.reg_window\[411\] final_design.cpu.reg_window\[443\] net960
+ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07730__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09343_ net474 _04098_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__or2_2
X_06555_ net752 _01505_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout241_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout339_A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09274_ net85 _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__or2_2
XFILLER_0_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06486_ final_design.reqhand.instruction\[19\] final_design.data_from_mem\[19\] net984
+ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__mux2_8
XFILLER_0_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06733__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14194__1263 vssd1 vssd1 vccd1 vccd1 _14194__1263/HI net1263 sky130_fd_sc_hd__conb_1
X_08225_ final_design.cpu.reg_window\[203\] final_design.cpu.reg_window\[235\] net856
+ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout506_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1248_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09588__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08156_ final_design.cpu.reg_window\[271\] final_design.cpu.reg_window\[303\] net827
+ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11395__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07107_ net896 _02051_ _02057_ _02044_ _02045_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__a32oi_4
XANTENNA__07063__A1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11934__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07685__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08087_ _01750_ _02896_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07038_ final_design.cpu.reg_window\[590\] final_design.cpu.reg_window\[622\] net935
+ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__mux2_1
XANTENNA__11147__A0 final_design.reqhand.data_from_UART\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14012__RESET_B net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08563__A1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ net627 _03921_ _03924_ _03655_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__B2 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11427__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07206__A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10951_ _05677_ _05678_ _05651_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_35_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13670_ clknet_leaf_170_clk _00901_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[658\]
+ sky130_fd_sc_hd__dfrtp_1
X_10882_ _05611_ _05612_ _05590_ _05593_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07640__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12621_ net1443 final_design.reqhand.data_from_UART\[7\] _05080_ vssd1 vssd1 vccd1
+ vccd1 _01314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _06215_ net359 net326 net1913 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__a22o_1
XANTENNA__11622__A1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10286__B net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ net2249 net229 net525 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12947__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12483_ _06143_ net343 net331 net2166 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14222_ final_design.h_out vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
X_11434_ net1811 net190 net313 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__mux2_1
XANTENNA__06780__A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09043__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11386__B1 _05947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11925__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14153_ clknet_leaf_78_clk _01327_ net1247 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11365_ net435 net589 _06053_ net317 net1791 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_100_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13104_ clknet_leaf_108_clk _00335_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[92\]
+ sky130_fd_sc_hd__dfrtp_1
X_10316_ net1550 net1022 net999 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1
+ vccd1 _00073_ sky130_fd_sc_hd__a22o_1
XANTENNA__06801__A1 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14084_ clknet_leaf_71_clk _01281_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11296_ _01881_ net649 _05991_ _05992_ net661 vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__a221o_1
X_13035_ clknet_leaf_14_clk _00266_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10247_ final_design.uart.BAUD_counter\[17\] final_design.uart.BAUD_counter\[16\]
+ _05114_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__and3_1
Xfanout1120 net1121 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12350__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1131 net1132 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_4
Xfanout1142 net1144 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__clkbuf_4
X_10178_ final_design.uart.BAUD_counter\[17\] final_design.uart.BAUD_counter\[16\]
+ final_design.uart.BAUD_counter\[19\] final_design.uart.BAUD_counter\[18\] vssd1
+ vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__or4_1
Xfanout1153 net1156 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08500__A _02330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1164 net100 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_4
XANTENNA__10361__B2 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1175 net1177 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__clkbuf_4
Xfanout1186 net1188 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06660__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1197 net1217 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08306__A1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_167_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_167_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13937_ clknet_leaf_91_clk _01168_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[925\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13868_ clknet_leaf_121_clk _01099_ net1197 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[856\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11861__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12819_ net1373 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11580__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12168__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13799_ clknet_leaf_16_clk _01030_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[787\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10416__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09282__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09985__B _04898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08010_ _02948_ _02949_ _02960_ net893 vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__a22o_4
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08381__S net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10924__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold603 final_design.cpu.reg_window\[183\] vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold614 final_design.cpu.reg_window\[487\] vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06479__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold625 final_design.cpu.reg_window\[780\] vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 final_design.cpu.reg_window\[869\] vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold647 final_design.cpu.reg_window\[878\] vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 final_design.cpu.reg_window\[578\] vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09961_ _04871_ _04876_ _04878_ net733 vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__a211o_2
Xhold669 final_design.cpu.reg_window\[553\] vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09417__S0 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08912_ _01692_ _02467_ net627 vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09892_ _02325_ net488 net444 vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12341__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09506__A _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ final_design.CPU_instr_adr\[19\] final_design.CPU_instr_adr\[18\] _03793_
+ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__and3_1
XANTENNA__06556__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout191_A _06038_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10352__B2 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout289_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ _03698_ _03724_ _03697_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07725_ final_design.cpu.reg_window\[282\] final_design.cpu.reg_window\[314\] net873
+ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_158_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_158_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11301__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07656_ net612 _02602_ _02577_ _01566_ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11490__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06607_ _01554_ _01555_ _01556_ _01557_ net786 net803 vssd1 vssd1 vccd1 vccd1 _01558_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07587_ _02534_ _02535_ _02536_ _02537_ net687 net708 vssd1 vssd1 vccd1 vccd1 _02538_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10407__A2 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09326_ _04056_ _04243_ _04244_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__o21a_1
X_06538_ _01456_ _01465_ _01474_ _01480_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__or4_4
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09257_ _04175_ net452 _04174_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__and3b_1
XFILLER_0_91_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06469_ final_design.reqhand.instruction\[15\] final_design.data_from_mem\[15\] net985
+ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout509_X net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08208_ net726 _03158_ net889 vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_170_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08291__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09188_ net493 _04055_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__nor2_2
XFILLER_0_161_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08139_ final_design.cpu.reg_window\[845\] final_design.cpu.reg_window\[877\] net834
+ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11011__A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _04805_ net665 _05843_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a211oi_4
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ final_design.vga.h_current_state\[0\] final_design.vga.h_current_state\[1\]
+ _05015_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11081_ net91 net1058 vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12332__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07635__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ _02836_ _04162_ _04158_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__or3b_1
XANTENNA__11665__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09135__B _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12096__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11983_ _06185_ net288 net406 net2097 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_149_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_149_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13722_ clknet_leaf_160_clk _00953_ net1105 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[710\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10934_ _01386_ _05649_ _05658_ _05661_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__nor4_1
XANTENNA__09422__Y _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07370__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13653_ clknet_leaf_53_clk _00884_ net1159 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[641\]
+ sky130_fd_sc_hd__dfrtp_1
X_10865_ net974 _05596_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__or2_1
X_12604_ net1411 net1010 net996 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1
+ vccd1 _01297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12399__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13584_ clknet_leaf_104_clk _00815_ net1204 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[572\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10796_ net76 _05511_ _05530_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12535_ _06198_ net353 net325 net1868 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12466_ _06126_ net350 net332 net2272 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__a22o_1
XANTENNA__06714__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14205_ net1274 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11417_ net1748 net244 net311 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__mux2_1
XANTENNA__09567__A3 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12397_ net564 _06268_ net341 net2089 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__a22o_1
X_14136_ clknet_leaf_77_clk final_design.vga.h_next_count\[5\] net1252 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[5\] sky130_fd_sc_hd__dfrtp_4
X_11348_ net657 net190 vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07983__C1 _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11856__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ clknet_leaf_46_clk net2553 net1147 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12451__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10760__A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ net653 _05977_ _05976_ net665 vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07545__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ clknet_leaf_164_clk _00249_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10334__B2 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06553__A3 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07750__A2 _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12087__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07510_ _01825_ _02460_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__or2_1
XANTENNA__07189__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08490_ final_design.cpu.reg_window\[963\] final_design.cpu.reg_window\[995\] net861
+ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07441_ final_design.reqhand.instruction\[8\] final_design.data_from_mem\[8\] net986
+ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08138__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10000__A _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07372_ _02319_ _02320_ _02321_ _02322_ net784 net793 vssd1 vssd1 vccd1 vccd1 _02323_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_91_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09111_ final_design.CPU_instr_adr\[0\] _02425_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10935__A _05662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12626__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11530__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09042_ net631 _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06624__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold400 final_design.reqhand.current_client\[0\] vssd1 vssd1 vccd1 vccd1 net1753
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 final_design.cpu.reg_window\[904\] vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout204_A _05989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold422 final_design.cpu.reg_window\[791\] vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 final_design.cpu.reg_window\[837\] vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12562__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold444 final_design.cpu.reg_window\[478\] vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold455 final_design.cpu.reg_window\[645\] vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold466 final_design.cpu.reg_window\[512\] vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold477 final_design.cpu.reg_window\[883\] vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold488 final_design.cpu.reg_window\[542\] vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout902 net903 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_4
X_09944_ _04861_ _04862_ _04858_ _04860_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__a2bb2o_2
Xfanout913 net917 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__clkbuf_4
Xhold499 final_design.cpu.reg_window\[233\] vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1113_A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08518__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout924 net933 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_4
Xfanout935 net936 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__buf_2
Xfanout946 net948 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ net536 net534 net455 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__mux2_1
Xfanout957 net965 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_4
Xfanout968 net970 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1100 final_design.cpu.reg_window\[317\] vssd1 vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10325__B2 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout573_A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 _04035_ vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__clkbuf_4
Xhold1111 final_design.cpu.reg_window\[564\] vssd1 vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 final_design.uart.working_data\[6\] vssd1 vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ final_design.CPU_instr_adr\[29\] _01539_ _03776_ vssd1 vssd1 vccd1 vccd1
+ _03777_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1133 final_design.cpu.reg_window\[651\] vssd1 vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1144 final_design.cpu.reg_window\[305\] vssd1 vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 final_design.cpu.reg_window\[307\] vssd1 vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 final_design.cpu.reg_window\[982\] vssd1 vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12078__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08757_ _03706_ _03707_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__nor2_1
Xhold1177 final_design.cpu.reg_window\[296\] vssd1 vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout740_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1188 final_design.cpu.reg_window\[292\] vssd1 vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1199 final_design.uart.BAUD_counter\[31\] vssd1 vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout838_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07708_ final_design.cpu.reg_window\[667\] final_design.cpu.reg_window\[699\] net879
+ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
X_08688_ net623 _03550_ _02419_ _02423_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_120_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06927__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ final_design.cpu.reg_window\[860\] final_design.cpu.reg_window\[892\] net874
+ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07978__X _02929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ _05368_ _05390_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11589__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09309_ _04091_ _04227_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__and2_1
X_10581_ _05326_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__inv_2
XANTENNA__11440__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12320_ net1775 net193 net364 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10564__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12251_ net587 _06180_ net515 net374 net1735 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11202_ _04903_ net659 net599 _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__o211a_2
XANTENNA__12553__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ net1730 net201 net380 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__mux2_1
XANTENNA__11761__A0 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ _05840_ _05846_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__or2_4
XFILLER_0_102_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07365__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ net1067 _05785_ _05786_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10316__B2 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _04220_ _04693_ _04932_ _04933_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_48_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08368__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11966_ _06168_ net282 net404 net2086 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ _05624_ _05646_ _05645_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__a21oi_1
X_13705_ clknet_leaf_95_clk _00936_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[693\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11897_ net212 net2100 net274 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13636_ clknet_leaf_98_clk _00867_ net1256 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[624\]
+ sky130_fd_sc_hd__dfrtp_1
X_10848_ _05578_ _05579_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14115__RESET_B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07248__A1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11044__A2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13567_ clknet_leaf_134_clk _00798_ net1167 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[555\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12446__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10779_ _05487_ _05489_ _05513_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__or3b_1
XFILLER_0_125_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09966__D _04884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12518_ _06180_ net356 net329 net1859 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13498_ clknet_leaf_163_clk _00729_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[486\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12449_ net2048 net204 net336 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11201__C1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12544__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14119_ clknet_leaf_76_clk final_design.vga.h_next_state\[1\] net1254 vssd1 vssd1
+ vccd1 vccd1 final_design.vga.h_current_state\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_35_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12181__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_2
X_07990_ final_design.cpu.reg_window\[400\] final_design.cpu.reg_window\[432\] net887
+ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__mux2_1
XANTENNA__13068__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06941_ final_design.cpu.reg_window\[209\] final_design.cpu.reg_window\[241\] net910
+ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09660_ _04362_ _04363_ net481 vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__o21ai_2
X_06872_ _01504_ _01822_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__nand2_2
XANTENNA__08895__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08611_ net535 _03386_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09591_ net736 _04482_ _04502_ _04508_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_141_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08542_ _03489_ _03490_ _03491_ _03492_ net689 net708 vssd1 vssd1 vccd1 vccd1 _03493_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_173_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11283__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ _03420_ _03422_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07424_ net770 _02374_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__or2_1
XFILLER_0_174_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12232__A1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07355_ final_design.cpu.reg_window\[67\] final_design.cpu.reg_window\[99\] net945
+ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07286_ _02233_ _02234_ _02235_ _02236_ net777 net797 vssd1 vssd1 vccd1 vccd1 _02237_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_171_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09025_ final_design.CPU_instr_adr\[12\] _03789_ vssd1 vssd1 vccd1 vccd1 _03957_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12535__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09936__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold230 net127 vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 final_design.VGA_data_control.ready_data\[14\] vssd1 vssd1 vccd1 vccd1 net1594
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout690_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 final_design.cpu.reg_window\[714\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 final_design.cpu.reg_window\[244\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold274 final_design.cpu.reg_window\[835\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 final_design.cpu.reg_window\[163\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold296 final_design.cpu.reg_window\[681\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 net716 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__buf_4
Xfanout721 net722 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__buf_4
XANTENNA__07185__S net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout732 _01688_ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_165_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12299__A1 _05875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09927_ _04843_ _04845_ _04831_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_165_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout743 net745 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__clkbuf_4
Xfanout754 net757 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__buf_6
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout955_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout765 _01427_ vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__buf_2
Xfanout776 net782 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_2
Xfanout787 net790 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_4
X_09858_ _03294_ net447 _04775_ _04776_ net263 vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__o2111ai_1
XANTENNA__09703__A3 _04579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout798 net807 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_4
X_08809_ final_design.CPU_instr_adr\[21\] _01788_ vssd1 vssd1 vccd1 vccd1 _03760_
+ sky130_fd_sc_hd__nand2_1
X_09789_ _04219_ _04343_ _04221_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a21o_1
XANTENNA__11435__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11820_ net218 net2043 net267 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11751_ net206 net2468 net416 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08675__B1 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10702_ _05438_ _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11682_ net425 net568 _06199_ net295 net1630 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__a32o_1
XFILLER_0_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13421_ clknet_leaf_140_clk _00652_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[409\]
+ sky130_fd_sc_hd__dfrtp_1
X_10633_ _05354_ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12223__A1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06772__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08978__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13352_ clknet_leaf_119_clk _00583_ net1199 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[340\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input84_A memory_size[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10564_ _04724_ net254 vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10785__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10785__B2 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11982__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ net1739 net237 net364 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13283_ clknet_leaf_4_clk _00514_ net1096 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[271\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07650__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10495_ _05234_ _05242_ _05243_ net58 vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_20_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12234_ net584 _06164_ net514 net374 net1803 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__a32o_1
XANTENNA__12526__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11734__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12165_ net2347 net229 net381 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07095__S net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11116_ final_design.uart.bits_received\[2\] _05832_ vssd1 vssd1 vccd1 vccd1 _05834_
+ sky130_fd_sc_hd__xnor2_1
X_12096_ net1886 net229 net389 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11047_ net978 _05770_ _05768_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_30_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07823__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12998_ net1340 _00229_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07013__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12462__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ _06150_ net289 net410 net1771 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_71_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10473__A0 final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12176__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12214__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ clknet_leaf_36_clk _00850_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[607\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10485__A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07140_ _02078_ _02079_ _02090_ net899 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_43_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11973__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07071_ final_design.cpu.reg_window\[973\] final_design.cpu.reg_window\[1005\] net915
+ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12517__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09615__B1_N _04231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09394__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07973_ final_design.cpu.reg_window\[657\] final_design.cpu.reg_window\[689\] net827
+ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__mux2_1
X_09712_ _04626_ _04630_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_143_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06924_ final_design.cpu.reg_window\[658\] final_design.cpu.reg_window\[690\] net901
+ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__mux2_1
X_09643_ net488 _04559_ _04560_ _04224_ _04092_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__a221o_1
X_06855_ final_design.cpu.reg_window\[916\] final_design.cpu.reg_window\[948\] net949
+ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout271_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout369_A net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09574_ _04492_ _04488_ net319 _04067_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__o2bb2a_1
X_06786_ net767 _01736_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__nor2_1
XANTENNA__14037__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08525_ final_design.cpu.reg_window\[642\] final_design.cpu.reg_window\[674\] net867
+ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12453__A1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout536_A _02239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ final_design.cpu.reg_window\[900\] final_design.cpu.reg_window\[932\] net859
+ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07407_ final_design.data_from_mem\[9\] net981 _02357_ vssd1 vssd1 vccd1 vccd1 _02358_
+ sky130_fd_sc_hd__o21a_2
XANTENNA__12205__A1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08387_ _03334_ _03335_ _03336_ _03337_ net685 net706 vssd1 vssd1 vccd1 vccd1 _03338_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout703_A _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_X net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07338_ final_design.cpu.reg_window\[644\] final_design.cpu.reg_window\[676\] net939
+ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11964__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07269_ _02216_ _02217_ _02218_ _02219_ net777 net797 vssd1 vssd1 vccd1 vccd1 _02220_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ net627 _03938_ net257 vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12508__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10280_ _05138_ net810 _05137_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_167_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11716__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09385__A1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_133_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 _02126_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__buf_2
Xfanout551 _01850_ vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_4
X_13970_ clknet_leaf_40_clk _01201_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[958\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout573 net574 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_4
Xfanout584 net585 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12769__B net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_4
XANTENNA__09424__A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ clknet_leaf_10_clk _00159_ net1092 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11673__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12692__A1 _05008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_148_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ clknet_leaf_86_clk _00090_ net1248 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11803_ net2493 net414 net289 _06046_ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__a22o_1
XANTENNA__12444__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11247__A2 _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11734_ net577 net422 _06225_ net296 net1782 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__a32o_1
XFILLER_0_139_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11665_ net178 net639 vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_25_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10616_ net1066 _05356_ net1014 final_design.CPU_instr_adr\[8\] vssd1 vssd1 vccd1
+ vccd1 _05360_ sky130_fd_sc_hd__o2bb2a_1
X_13404_ clknet_leaf_147_clk _00635_ net1127 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[392\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input87_X net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11596_ net180 net645 vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__and2_1
XANTENNA__10302__S0 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11955__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13335_ clknet_leaf_141_clk _00566_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[323\]
+ sky130_fd_sc_hd__dfrtp_1
X_10547_ _05273_ _05292_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13342__RESET_B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13266_ clknet_leaf_38_clk _00497_ net1136 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[254\]
+ sky130_fd_sc_hd__dfrtp_1
X_10478_ net47 _05223_ _05225_ _05227_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__and4_1
XFILLER_0_122_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12217_ net587 _06145_ net516 net378 net1680 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__a32o_1
X_13197_ clknet_leaf_140_clk _00428_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[185\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09915__A3 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11183__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ net201 net2484 net384 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ net568 _05990_ net505 net392 net1901 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12132__A0 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12683__B2 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10694__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ final_design.cpu.reg_window\[667\] final_design.cpu.reg_window\[699\] net958
+ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__mux2_1
XANTENNA__14130__RESET_B net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12435__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06571_ net765 _01515_ net757 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_47_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08310_ net619 _03257_ _03258_ net539 vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09290_ _02639_ net444 net440 _02638_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__o22a_1
XANTENNA__08384__S net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08241_ _03179_ _03180_ _03191_ net892 vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_118_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12199__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08172_ final_design.cpu.reg_window\[719\] final_design.cpu.reg_window\[751\] net824
+ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09603__A2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11946__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07123_ final_design.cpu.reg_window\[11\] final_design.cpu.reg_window\[43\] net937
+ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__mux2_1
XANTENNA__11598__X _06155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07054_ final_design.cpu.reg_window\[461\] final_design.cpu.reg_window\[493\] net914
+ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__clkbuf_4
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
XANTENNA__11174__A1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1026_A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout486_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ final_design.cpu.reg_window\[273\] final_design.cpu.reg_window\[305\] net836
+ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06907_ final_design.cpu.reg_window\[274\] final_design.cpu.reg_window\[306\] net903
+ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07225__S0 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07887_ _02800_ _02801_ _02833_ _02835_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06838_ _01785_ _01788_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__nor2_1
X_09626_ _02868_ _04544_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_108_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09557_ _04474_ _04475_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11229__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06769_ final_design.data_from_mem\[23\] net981 _01719_ vssd1 vssd1 vccd1 vccd1 _01720_
+ sky130_fd_sc_hd__o21a_2
XANTENNA_fanout820_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_X net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout918_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08508_ final_design.cpu.reg_window\[258\] final_design.cpu.reg_window\[290\] net866
+ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__mux2_1
XANTENNA__10437__B1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09488_ net478 _04406_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__nor2_1
XANTENNA__08294__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08439_ _03387_ _03389_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11014__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08763__B1_N final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11450_ net227 net647 vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__and2_1
XANTENNA__11937__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10401_ net1430 net1040 _05183_ net246 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11381_ net657 net183 vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__and2_2
X_13120_ clknet_leaf_36_clk _00351_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_12_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ net1585 net1023 net1000 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1
+ vccd1 _00089_ sky130_fd_sc_hd__a22o_1
XANTENNA__08323__A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13051_ clknet_leaf_156_clk _00282_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_10263_ final_design.uart.BAUD_counter\[23\] final_design.uart.BAUD_counter\[22\]
+ _05124_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__and3_1
X_12002_ _06204_ net287 net401 net1601 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__a22o_1
XANTENNA__12362__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input47_A mem_adr_start[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ final_design.uart.BAUD_counter\[1\] final_design.uart.BAUD_counter\[0\] vssd1
+ vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__or2_1
XANTENNA__10912__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10912__B2 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout370 net371 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout381 net383 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_6
Xfanout392 net393 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_8
X_13953_ clknet_leaf_158_clk _01184_ net1113 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[941\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12665__B2 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12904_ clknet_leaf_11_clk _00142_ net1092 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
X_13884_ clknet_leaf_147_clk _01115_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[872\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12835_ clknet_leaf_72_clk _00073_ net1245 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10428__B1 _05197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12766_ _06383_ _06396_ _06397_ _06400_ _06401_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__a311o_1
XANTENNA__10979__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10979__B2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11717_ net192 net634 vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__and2_1
X_12697_ final_design.VGA_data_control.v_count\[8\] final_design.VGA_data_control.v_count\[5\]
+ _01398_ _06336_ final_design.VGA_data_control.v_count\[7\] vssd1 vssd1 vccd1 vccd1
+ _06338_ sky130_fd_sc_hd__a32o_1
XANTENNA__11640__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08217__B net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11648_ net595 net424 _06181_ net302 net1643 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11928__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput34 en vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
XANTENNA__09141__S0 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput45 mem_adr_start[18] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12454__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11579_ net434 net586 _06145_ net305 net2008 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__a32o_1
Xinput56 mem_adr_start[28] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput67 mem_adr_start[9] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__buf_1
XANTENNA__11211__X _05918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold807 final_design.cpu.reg_window\[182\] vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
Xinput78 memory_size[19] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07548__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput89 memory_size[29] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_4
Xhold818 final_design.cpu.reg_window\[802\] vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ clknet_leaf_168_clk _00549_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[306\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11578__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold829 final_design.cpu.reg_window\[536\] vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12026__Y _06261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13249_ clknet_leaf_162_clk _00480_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[237\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11156__A1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12353__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10903__A1 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07810_ _02757_ _02758_ _02759_ _02760_ net691 net702 vssd1 vssd1 vccd1 vccd1 _02761_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11594__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08790_ _03685_ _03686_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__nand2_1
XANTENNA__08379__S net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08309__C1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ final_design.cpu.reg_window\[730\] final_design.cpu.reg_window\[762\] net872
+ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07672_ net719 _02616_ net732 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__o21a_1
X_09411_ _04158_ _04163_ _02837_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06623_ final_design.cpu.reg_window\[475\] final_design.cpu.reg_window\[507\] net961
+ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_17_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11533__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ net473 _04260_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_138_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06554_ final_design.reqhand.instruction\[30\] final_design.data_from_mem\[30\] net983
+ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__mux2_2
XANTENNA__08088__A1 _01718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06627__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09273_ net83 net84 _04191_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__or3_1
X_06485_ net769 _01435_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_62_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08224_ final_design.cpu.reg_window\[11\] final_design.cpu.reg_window\[43\] net856
+ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11919__B1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08155_ final_design.cpu.reg_window\[335\] final_design.cpu.reg_window\[367\] net827
+ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout401_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12364__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_151_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09884__D _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1143_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07106_ net769 _02056_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__or2_1
XANTENNA__11488__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08086_ _03035_ _03036_ _02901_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07037_ net760 _01987_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11147__A1 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_X net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12344__B1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08012__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__X _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout770_A _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__A2 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08289__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ net630 _03923_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__or2_1
X_07939_ final_design.cpu.reg_window\[598\] final_design.cpu.reg_window\[630\] net819
+ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__mux2_1
XANTENNA__12647__B2 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10950_ net84 net1060 vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__or2_1
XANTENNA__07206__B _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09609_ _04513_ _04527_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_27_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10881_ net81 _05589_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_158_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11870__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12620_ final_design.uart.working_data\[7\] net1414 _05080_ vssd1 vssd1 vccd1 vccd1
+ _01313_ sky130_fd_sc_hd__mux2_1
XANTENNA__09421__B _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12551_ _06214_ net355 net325 net2296 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11622__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10286__C _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11502_ net1781 net230 net526 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12482_ _06142_ net352 net332 net2135 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14221_ net1290 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
X_11433_ net1774 net192 net312 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07368__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14152_ clknet_leaf_80_clk _01326_ net1251 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11364_ net656 net186 vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__and2_1
XANTENNA__12987__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10315_ net1567 net1022 net999 final_design.data_from_mem\[0\] vssd1 vssd1 vccd1
+ vccd1 _00072_ sky130_fd_sc_hd__a22o_1
X_13103_ clknet_leaf_92_clk _00334_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[91\]
+ sky130_fd_sc_hd__dfrtp_1
X_14083_ clknet_leaf_71_clk _01280_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11295_ net743 _03909_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__nand2_1
XANTENNA__08988__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12335__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ clknet_leaf_1_clk _00265_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10246_ final_design.uart.BAUD_counter\[15\] final_design.uart.BAUD_counter\[16\]
+ _05113_ final_design.uart.BAUD_counter\[17\] vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__a31o_1
Xfanout1110 net1111 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__buf_2
Xfanout1121 net1128 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09751__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1132 net1137 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_2
X_10177_ final_design.uart.BAUD_counter\[21\] final_design.uart.BAUD_counter\[20\]
+ final_design.uart.BAUD_counter\[23\] final_design.uart.BAUD_counter\[22\] vssd1
+ vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__or4_1
XANTENNA__08199__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1143 net1144 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__clkbuf_4
Xfanout1154 net1156 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__clkbuf_4
Xfanout1165 net1168 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__clkbuf_4
Xfanout1176 net1177 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06660__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1187 net1188 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__clkbuf_4
Xfanout1198 net1200 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13936_ clknet_leaf_111_clk _01167_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[924\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11310__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07831__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09612__A _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10758__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12449__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867_ clknet_leaf_19_clk _01098_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[855\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11861__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12818_ net1358 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11580__C net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08228__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13798_ clknet_leaf_168_clk _01029_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[786\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11074__B1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12749_ _06381_ _06383_ _06384_ _06387_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09282__A3 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09019__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10493__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12184__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07278__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold604 final_design.cpu.reg_window\[241\] vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 final_design.cpu.reg_window\[551\] vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06479__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold626 final_design.cpu.reg_window\[468\] vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold637 final_design.cpu.reg_window\[189\] vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold648 final_design.cpu.reg_window\[985\] vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 final_design.cpu.reg_window\[65\] vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09960_ _04871_ _04876_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08911_ final_design.CPU_instr_adr\[25\] net1029 _03851_ _03855_ vssd1 vssd1 vccd1
+ vccd1 _00236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09891_ _04147_ _04809_ net450 vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a21o_1
XANTENNA__11528__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10888__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ final_design.CPU_instr_adr\[17\] _03792_ vssd1 vssd1 vccd1 vccd1 _03793_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06556__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10352__A2 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08773_ _03701_ _03722_ _03700_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_109_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12629__B2 final_design.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout184_A _06060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07724_ final_design.cpu.reg_window\[346\] final_design.cpu.reg_window\[378\] net872
+ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__mux2_1
XANTENNA__11301__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07741__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08702__C1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07655_ _01567_ _02604_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07600__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1093_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06606_ final_design.cpu.reg_window\[924\] final_design.cpu.reg_window\[956\] net954
+ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout449_A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07586_ final_design.cpu.reg_window\[927\] final_design.cpu.reg_window\[959\] net841
+ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09325_ net265 _04217_ _04230_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__and3_1
X_06537_ _01456_ _01465_ _01473_ _01481_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_153_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout237_X net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout616_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09256_ _02638_ _04173_ _02545_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__a21boi_1
X_06468_ final_design.data_from_mem\[17\] net982 _01417_ vssd1 vssd1 vccd1 vccd1 _01419_
+ sky130_fd_sc_hd__o21ai_4
XANTENNA_clkbuf_4_10__f_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08207_ _03154_ _03155_ _03156_ _03157_ net688 net701 vssd1 vssd1 vccd1 vccd1 _03158_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09187_ _03519_ _04104_ _04105_ _04098_ net474 vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_90_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__A1 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1146_X net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07188__S net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08138_ _03085_ _03086_ _03087_ _03088_ net685 net706 vssd1 vssd1 vccd1 vccd1 _03089_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout985_A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08784__A2 _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08069_ _03016_ _03017_ _03018_ _03019_ net682 net699 vssd1 vssd1 vccd1 vccd1 _03020_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10100_ _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__inv_2
X_11080_ net1058 net91 vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11438__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ net322 _04949_ _04948_ _04947_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__o211a_1
XANTENNA__08536__A2 _03481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14111__Q final_design.reqhand.data_from_UART\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11982_ _06184_ net290 net406 net1569 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11681__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ clknet_leaf_165_clk _00952_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[709\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10933_ _05649_ _05658_ _05661_ _01386_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__o31a_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09151__B _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ net968 _05585_ _05595_ net972 vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__o22a_1
X_13652_ clknet_leaf_104_clk _00883_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[640\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12603_ net1387 net1010 net996 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1
+ vccd1 _01296_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _05528_ _05529_ _05511_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_54_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13583_ clknet_leaf_92_clk _00814_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[571\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11901__S net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12534_ _06197_ net354 net325 net1897 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__a22o_1
XANTENNA__08482__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12465_ net680 net645 _06268_ net334 net2233 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__a32o_1
XANTENNA__11359__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12556__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14204_ net1273 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11416_ net1942 net237 net311 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12396_ net563 net507 vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__nand2_1
XANTENNA__10031__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14135_ clknet_leaf_75_clk final_design.vga.h_next_count\[4\] net1253 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[4\] sky130_fd_sc_hd__dfrtp_1
X_11347_ _06034_ _06036_ _06037_ net599 vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__o211a_4
XFILLER_0_120_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07826__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09607__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14066_ clknet_leaf_46_clk _00029_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11278_ final_design.data_from_mem\[16\] _05177_ _05912_ _05917_ vssd1 vssd1 vccd1
+ vccd1 _05977_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06730__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11856__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ net2220 _05104_ _05106_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__a21oi_1
X_13017_ clknet_leaf_167_clk _00248_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07735__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11531__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07127__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 wb_manage.BUSY_O vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11872__A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06553__A4 _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10098__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09342__A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13919_ clknet_leaf_135_clk _01150_ net1167 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[907\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10488__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12179__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07440_ _01489_ net741 _01495_ net697 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a31o_1
XFILLER_0_159_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08138__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07371_ final_design.cpu.reg_window\[515\] final_design.cpu.reg_window\[547\] net942
+ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09110_ _04030_ final_design.CPU_instr_adr\[1\] _03812_ vssd1 vssd1 vccd1 vccd1 _00210_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11811__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09041_ _03730_ _03970_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12547__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold401 final_design.cpu.reg_window\[72\] vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12011__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07649__S0 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold412 final_design.cpu.reg_window\[194\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold423 final_design.cpu.reg_window\[924\] vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 final_design.cpu.reg_window\[576\] vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold445 final_design.cpu.reg_window\[853\] vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold456 final_design.cpu.reg_window\[964\] vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07736__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold467 final_design.cpu.reg_window\[912\] vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold478 final_design.cpu.reg_window\[902\] vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold489 final_design.cpu.reg_window\[409\] vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ _03390_ _03421_ _04149_ net450 vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__a31o_1
Xfanout903 net912 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_2
Xfanout914 net917 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout925 net933 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_4
Xfanout936 net966 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_74_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout399_A _06261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout947 net948 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10015__X _04934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ _04460_ _04465_ _04727_ _04461_ _04222_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_146_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout958 net965 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__clkbuf_4
Xfanout969 net970 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 final_design.cpu.reg_window\[614\] vssd1 vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1106_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1112 final_design.cpu.reg_window\[35\] vssd1 vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07037__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09804__X _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1123 final_design.reqhand.instruction\[2\] vssd1 vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ final_design.CPU_instr_adr\[28\] _01570_ _03775_ vssd1 vssd1 vccd1 vccd1
+ _03776_ sky130_fd_sc_hd__a21o_1
Xhold1134 final_design.cpu.reg_window\[130\] vssd1 vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1145 final_design.cpu.reg_window\[318\] vssd1 vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 final_design.cpu.reg_window\[944\] vssd1 vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 final_design.cpu.reg_window\[482\] vssd1 vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08756_ _01366_ _02297_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__and2_1
Xhold1178 final_design.cpu.reg_window\[260\] vssd1 vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1189 final_design.cpu.reg_window\[994\] vssd1 vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07707_ final_design.cpu.reg_window\[731\] final_design.cpu.reg_window\[763\] net881
+ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout733_A _01493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ _03456_ _03457_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_120_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ net728 _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout900_A _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07569_ _02516_ _02517_ _02518_ _02519_ net688 net709 vssd1 vssd1 vccd1 vccd1 _02520_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11589__A1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09308_ net530 net493 vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10580_ net64 _05324_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09239_ _02936_ _04135_ _04143_ _04157_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__or4_4
XFILLER_0_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12538__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_9__f_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12250_ net570 _06179_ net506 net372 net1629 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_118_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12002__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11201_ _05855_ _05906_ _05908_ net663 vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__a211o_1
XANTENNA__11957__A net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ net2177 net203 net380 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ _05840_ _05846_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__nor2_4
XFILLER_0_102_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold990 final_design.reqhand.instruction\[9\] vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11168__S net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11063_ final_design.CPU_instr_adr\[29\] net1054 net814 vssd1 vssd1 vccd1 vccd1 _05786_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__08914__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ net490 _04779_ _04341_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_4_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10800__S net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06786__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07234__X _02185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08368__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11965_ _06167_ net282 net404 net1624 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ clknet_leaf_117_clk _00935_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[692\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10916_ net49 _05620_ _05625_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_80_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11896_ net214 net2205 net276 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ clknet_leaf_1_clk _00866_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[623\]
+ sky130_fd_sc_hd__dfrtp_1
X_10847_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06725__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13566_ clknet_leaf_18_clk _00797_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[554\]
+ sky130_fd_sc_hd__dfrtp_1
X_10778_ _05487_ _05489_ _05513_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_171_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09101__S net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12517_ _06179_ net345 net327 net1935 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__a22o_1
X_13497_ clknet_leaf_165_clk _00728_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[485\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12529__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12448_ net1820 net221 net338 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12462__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12379_ net1945 net206 net270 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__mux2_1
X_14118_ clknet_leaf_76_clk final_design.vga.h_next_state\[0\] net1254 vssd1 vssd1
+ vccd1 vccd1 final_design.vga.h_current_state\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__11586__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06940_ final_design.cpu.reg_window\[17\] final_design.cpu.reg_window\[49\] net910
+ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__mux2_1
X_14049_ clknet_leaf_48_clk _00010_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11504__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06871_ net751 net674 _01819_ _01821_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08610_ _03455_ _03557_ _03560_ _03457_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__o31a_1
X_09590_ _04502_ _04508_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__nand2_2
XANTENNA__10489__Y _05239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07144__X _02095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11268__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08541_ final_design.cpu.reg_window\[385\] final_design.cpu.reg_window\[417\] net849
+ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__mux2_1
XANTENNA__11807__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08133__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08472_ _03420_ _03422_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__nor2_1
XANTENNA__12480__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09881__B1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07423_ _02370_ _02371_ _02372_ _02373_ net781 net799 vssd1 vssd1 vccd1 vccd1 _02374_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_92_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10491__A1 _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10491__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10946__A _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12787__18 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__inv_2
X_07354_ _02301_ _02302_ _02303_ _02304_ net784 net802 vssd1 vssd1 vccd1 vccd1 _02305_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07285_ final_design.cpu.reg_window\[646\] final_design.cpu.reg_window\[678\] net913
+ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout314_A _06092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09024_ net627 _03955_ _03954_ net256 vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08703__X _03654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold220 net164 vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12372__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold231 final_design.cpu.reg_window\[220\] vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1223_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold242 final_design.VGA_data_control.ready_data\[26\] vssd1 vssd1 vccd1 vccd1 net1595
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold253 final_design.cpu.reg_window\[699\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 final_design.cpu.reg_window\[184\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 final_design.cpu.reg_window\[540\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold286 final_design.cpu.reg_window\[62\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout700 net701 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_2
XANTENNA_fanout683_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold297 net125 vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 net714 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout722 net723 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_4
X_09926_ _04124_ _04718_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_165_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout733 _01493_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_4
Xfanout744 net745 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_2
Xfanout755 net757 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_4
Xfanout777 net778 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_8
X_09857_ _03292_ net443 net439 _03291_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__o22a_1
XANTENNA__07175__A1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout788 net789 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_4
Xfanout799 net801 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__buf_4
XANTENNA_fanout948_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08911__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ _03757_ _03758_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__and2_1
XANTENNA__08297__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09788_ _03358_ _04705_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__xnor2_1
X_08739_ final_design.CPU_instr_adr\[10\] _02128_ vssd1 vssd1 vccd1 vccd1 _03690_
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08675__A1 _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11750_ net208 net1988 net416 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__mux2_1
XANTENNA__09872__B1 _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ _05404_ _05439_ _05440_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_166_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11681_ net224 net634 vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__and2_1
XANTENNA__11451__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13420_ clknet_leaf_119_clk _00651_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[408\]
+ sky130_fd_sc_hd__dfrtp_1
X_10632_ _05372_ _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10563_ _05268_ _05305_ _05307_ _05302_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13351_ clknet_leaf_16_clk _00582_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[339\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_950 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14192__1262 vssd1 vssd1 vccd1 vccd1 _14192__1262/HI net1262 sky130_fd_sc_hd__conb_1
XFILLER_0_107_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12302_ net1806 net224 net364 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input77_A memory_size[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10494_ net58 _05234_ _05242_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__and4_1
X_13282_ clknet_leaf_21_clk _00513_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[270\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12233_ net585 _06163_ net517 net374 net1460 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__a32o_1
XANTENNA__08286__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ net1747 net231 net382 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__mux2_1
XANTENNA__08699__C _03649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ final_design.uart.bits_received\[1\] _05830_ _05831_ _05833_ vssd1 vssd1
+ vccd1 vccd1 _00206_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ net1787 net231 net390 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__mux2_1
XANTENNA__08038__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11046_ net971 _05767_ _05769_ net969 vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08000__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12997_ net1339 _00228_ net1159 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07469__A2 _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08666__A1 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ _06149_ net290 net410 net2082 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__a22o_1
XANTENNA__07013__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12457__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11879_ _06113_ net291 net522 net2062 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11214__X _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13618_ clknet_leaf_42_clk _00849_ net1150 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[606\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09091__A1 final_design.CPU_instr_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13549_ clknet_leaf_137_clk _00780_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[537\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07070_ final_design.cpu.reg_window\[781\] final_design.cpu.reg_window\[813\] net917
+ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12192__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07972_ final_design.cpu.reg_window\[721\] final_design.cpu.reg_window\[753\] net827
+ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09711_ _04628_ _04629_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__nor2_2
XANTENNA__11489__A0 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06923_ final_design.cpu.reg_window\[722\] final_design.cpu.reg_window\[754\] net901
+ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__mux2_1
X_09642_ net488 _04559_ _04560_ _04262_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__a22o_1
X_06854_ final_design.cpu.reg_window\[980\] final_design.cpu.reg_window\[1012\] net956
+ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06785_ _01732_ _01733_ _01734_ _01735_ net774 net795 vssd1 vssd1 vccd1 vccd1 _01736_
+ sky130_fd_sc_hd__mux4_1
X_09573_ net499 net486 _04491_ _04409_ _04101_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__o32a_1
XFILLER_0_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout264_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08524_ final_design.cpu.reg_window\[706\] final_design.cpu.reg_window\[738\] net865
+ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08201__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09530__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08455_ final_design.cpu.reg_window\[964\] final_design.cpu.reg_window\[996\] net858
+ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__mux2_1
XANTENNA__12367__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10676__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout431_A _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1173_A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07406_ final_design.reqhand.instruction\[9\] net983 vssd1 vssd1 vccd1 vccd1 _02357_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_163_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08386_ final_design.cpu.reg_window\[134\] final_design.cpu.reg_window\[166\] net831
+ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_978 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07337_ final_design.cpu.reg_window\[708\] final_design.cpu.reg_window\[740\] net939
+ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09529__X _04448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07268_ final_design.cpu.reg_window\[390\] final_design.cpu.reg_window\[422\] net914
+ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__mux2_1
XANTENNA__08580__S net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout898_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ _02451_ net627 _03937_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07199_ final_design.cpu.reg_window\[521\] final_design.cpu.reg_window\[553\] net923
+ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11177__C1 _05887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11300__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774__5 clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__inv_2
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout530 _02502_ vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_4
Xfanout541 net542 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_2
X_09909_ _04806_ _04807_ _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__and3_1
Xfanout552 _01815_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_2
Xfanout563 _06238_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_4
Xfanout574 net575 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout585 net597 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12920_ clknet_leaf_10_clk _00158_ net1092 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dfrtp_1
Xfanout596 net597 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_2
X_12851_ clknet_leaf_86_clk _00089_ net1248 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11802_ net2506 net414 net290 _06039_ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09711__Y _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11652__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10455__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11733_ net176 net635 vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__and2_1
XANTENNA__10586__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11664_ net437 net592 _06189_ net302 net1480 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__a32o_1
XFILLER_0_148_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13403_ clknet_leaf_153_clk _00634_ net1117 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[391\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10615_ net977 _05358_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11595_ net435 net589 _06153_ net305 net1591 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__a32o_1
XANTENNA__10302__S1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13334_ clknet_leaf_128_clk _00565_ net1192 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[322\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10546_ _05273_ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08490__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ clknet_leaf_107_clk _00496_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[253\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_94_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10477_ _05223_ _05225_ _05227_ net47 vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12216_ net570 _06144_ net506 net376 net2037 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__a32o_1
X_13196_ clknet_leaf_123_clk _00427_ net1191 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[184\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12147_ net203 net2469 net384 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12078_ net594 _05981_ net518 net395 net1853 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__a32o_1
X_11029_ _05752_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__inv_2
XANTENNA__08431__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12683__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09902__X _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__A0 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06898__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06570_ net773 _01520_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_47_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12187__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08240_ _03185_ _03190_ net722 vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12199__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08171_ _03118_ _03119_ _03120_ _03121_ net683 net705 vssd1 vssd1 vccd1 vccd1 _03122_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_83_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07122_ final_design.cpu.reg_window\[75\] final_design.cpu.reg_window\[107\] net937
+ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06913__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07053_ final_design.cpu.reg_window\[269\] final_design.cpu.reg_window\[301\] net917
+ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__clkbuf_4
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_110_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_162_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1019_A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ final_design.cpu.reg_window\[337\] final_design.cpu.reg_window\[369\] net836
+ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout381_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06868__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12123__A1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06906_ final_design.cpu.reg_window\[338\] final_design.cpu.reg_window\[370\] net905
+ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__mux2_1
X_07886_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__inv_2
XANTENNA__07225__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11331__C1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14191__1261 vssd1 vssd1 vccd1 vccd1 _14191__1261/HI net1261 sky130_fd_sc_hd__conb_1
X_09625_ _02900_ _04353_ _03038_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__a21oi_1
X_06837_ net749 net690 _01504_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__o21ai_4
XANTENNA__11882__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout267_X net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout646_A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06984__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09556_ net76 _04187_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__xor2_1
X_06768_ final_design.reqhand.instruction\[23\] net984 vssd1 vssd1 vccd1 vccd1 _01719_
+ sky130_fd_sc_hd__or2_1
XANTENNA__08575__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12426__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09260__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08507_ final_design.cpu.reg_window\[322\] final_design.cpu.reg_window\[354\] net866
+ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__mux2_1
XANTENNA__12097__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11634__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout813_A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06699_ net762 _01649_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__or2_1
X_09487_ _04404_ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08438_ net611 _03384_ _03360_ net535 vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_156_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08369_ _03314_ _03319_ net724 vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07919__S net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10400_ net528 _05181_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__nor2_1
X_11380_ _06063_ _06065_ _06066_ net599 vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__o211a_2
XFILLER_0_117_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07161__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10331_ net1487 net1023 net1000 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1
+ vccd1 _00088_ sky130_fd_sc_hd__a22o_1
XANTENNA__13822__RESET_B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10262_ final_design.uart.BAUD_counter\[21\] final_design.uart.BAUD_counter\[22\]
+ _05123_ final_design.uart.BAUD_counter\[23\] vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__a31o_1
X_13050_ clknet_leaf_163_clk _00281_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12001_ _06203_ net284 net401 net1953 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__a22o_1
X_10193_ final_design.uart.bits_received\[0\] final_design.uart.bits_received\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout360 net361 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_8
Xfanout371 _06274_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_8
Xfanout382 net383 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_8
X_13952_ clknet_leaf_38_clk _01183_ net1136 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[940\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout393 _06263_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12665__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12903_ clknet_leaf_100_clk _00141_ net1187 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_2
X_13883_ clknet_leaf_154_clk _01114_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[871\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11904__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12834_ clknet_leaf_72_clk _00072_ net1245 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12417__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10428__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12765_ final_design.VGA_adr\[7\] net808 vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11205__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11716_ net425 net567 _06216_ net295 net2057 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__a32o_1
XFILLER_0_84_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12696_ final_design.VGA_data_control.v_count\[8\] _01398_ vssd1 vssd1 vccd1 vccd1
+ _06337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11647_ net600 _06016_ net641 vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_42_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_1
XFILLER_0_24_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07829__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput35 gpio_in[5] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09141__S1 _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput46 mem_adr_start[19] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_1
X_11578_ net198 net644 vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__and2_1
Xinput57 mem_adr_start[29] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_1
Xinput68 memory_size[0] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06804__B1 _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold808 final_design.cpu.reg_window\[498\] vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13317_ clknet_leaf_150_clk _00548_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[305\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput79 memory_size[1] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_1
X_10529_ net1072 _03784_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold819 final_design.cpu.reg_window\[247\] vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13248_ clknet_leaf_35_clk _00479_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[236\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11875__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10364__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ clknet_leaf_157_clk _00410_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[167\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10903__A2 _05610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11594__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11086__S net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07780__B2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ _02687_ _02688_ _02689_ _02690_ net694 net713 vssd1 vssd1 vccd1 vccd1 _02691_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_165_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11313__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07671_ net726 _02621_ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__or2_1
XANTENNA__06966__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ _04289_ _04290_ _04327_ _04328_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__and4_1
XANTENNA__11814__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06622_ final_design.cpu.reg_window\[283\] final_design.cpu.reg_window\[315\] net961
+ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12408__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06553_ _01485_ _01489_ net741 _01495_ _01502_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__a41o_4
XANTENNA__11616__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ _04258_ _04259_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_138_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09285__A1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09272_ net82 _04190_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__or2_2
X_06484_ _01431_ _01432_ _01433_ _01434_ net779 net800 vssd1 vssd1 vccd1 vccd1 _01435_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_132_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07391__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08223_ final_design.cpu.reg_window\[75\] final_design.cpu.reg_window\[107\] net856
+ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11919__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout227_A _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07739__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08245__C1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ _01967_ net606 vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_151_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07105_ _02052_ _02053_ _02054_ _02055_ net779 net792 vssd1 vssd1 vccd1 vccd1 _02056_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12592__B2 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08085_ _01785_ _02799_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1136_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_147_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07036_ _01983_ _01984_ _01985_ _01986_ net780 net799 vssd1 vssd1 vccd1 vccd1 _01987_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout596_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__S net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08012__A2 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07220__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _03747_ _03922_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout763_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ final_design.cpu.reg_window\[662\] final_design.cpu.reg_window\[694\] net819
+ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11855__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07869_ final_design.cpu.reg_window\[980\] final_design.cpu.reg_window\[1012\] net868
+ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09608_ _04254_ _04514_ _04526_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_158_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10880_ _05609_ _05610_ _05589_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__o21bai_1
XANTENNA__14021__RESET_B net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11870__A3 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09539_ net556 net555 net554 net553 net454 net463 vssd1 vssd1 vccd1 vccd1 _04458_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_159_Left_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12550_ _06213_ net345 net323 net2291 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__a22o_1
XANTENNA__12280__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11501_ net527 vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ _06141_ net358 net333 net2509 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__a22o_1
XANTENNA__11312__X _06007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14220_ net1289 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_163_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11432_ net2103 net194 net311 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11679__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12127__Y _06266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12583__B2 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151_ clknet_leaf_80_clk _01325_ net1249 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11363_ _04528_ _05143_ net599 _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__o211a_2
XFILLER_0_132_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13102_ clknet_leaf_115_clk _00333_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_10314_ _05165_ net1022 vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14082_ clknet_leaf_71_clk _01279_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11294_ net667 _03906_ net739 vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_168_Left_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11695__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13033_ clknet_leaf_95_clk _00264_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10245_ net1810 _05114_ _05116_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10346__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1100 net1103 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07384__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1111 net1128 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__clkbuf_2
X_10176_ net1065 _05065_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__and2_2
Xfanout1122 net1124 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1133 net1137 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__clkbuf_4
Xfanout1144 net1145 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__buf_2
Xfanout1155 net1156 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__buf_2
Xfanout1166 net1168 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10104__A final_design.VGA_data_control.v_count\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1177 net1189 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__buf_2
Xfanout190 _06038_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_2
Xfanout1188 net1189 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__clkbuf_4
Xfanout1199 net1200 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_117_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13935_ clknet_leaf_89_clk _01166_ net1233 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[923\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11846__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload5_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13866_ clknet_leaf_165_clk _01097_ net1085 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[854\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11861__A3 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12817_ net1408 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_83_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13797_ clknet_leaf_151_clk _01028_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[785\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12748_ net967 _05058_ _06359_ _06372_ _06386_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__a41o_1
XANTENNA__12271__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10821__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10821__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12679_ final_design.VGA_data_control.ready_data\[27\] net1034 net989 final_design.data_from_mem\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_13_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11222__X _05928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12023__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14190__1260 vssd1 vssd1 vccd1 vccd1 _14190__1260/HI net1260 sky130_fd_sc_hd__conb_1
Xhold605 final_design.cpu.reg_window\[525\] vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10585__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold616 final_design.cpu.reg_window\[481\] vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold627 final_design.cpu.reg_window\[382\] vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold638 final_design.cpu.reg_window\[992\] vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 final_design.cpu.reg_window\[79\] vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08910_ net259 _03853_ net1029 vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10713__S net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10337__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09890_ _03638_ _04146_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__or2_1
XANTENNA__06699__A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08841_ final_design.CPU_instr_adr\[16\] final_design.CPU_instr_adr\[15\] _03791_
+ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08772_ _03702_ _03722_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__nand2_1
XANTENNA__09803__A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07723_ _01630_ net610 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__nand2_1
XANTENNA__10949__A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_A _06089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07654_ net626 _02602_ _02603_ _01566_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a211oi_1
XANTENNA__07600__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06605_ final_design.cpu.reg_window\[988\] final_design.cpu.reg_window\[1020\] net954
+ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07585_ final_design.cpu.reg_window\[991\] final_design.cpu.reg_window\[1023\] net845
+ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout344_A net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09324_ _04234_ _04242_ net495 vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__mux2_1
X_06536_ _01456_ _01465_ _01474_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__or3_4
XANTENNA__12262__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09255_ _02545_ _02637_ _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__or3b_1
X_06467_ final_design.data_from_mem\[17\] net981 _01417_ vssd1 vssd1 vccd1 vccd1 _01418_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout511_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12375__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout609_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13414__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ final_design.cpu.reg_window\[526\] final_design.cpu.reg_window\[558\] net853
+ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12014__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09186_ net562 net469 net456 vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_170_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08154__A _01967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08137_ final_design.cpu.reg_window\[653\] final_design.cpu.reg_window\[685\] net832
+ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__mux2_1
XANTENNA__09430__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1041_X net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08068_ final_design.cpu.reg_window\[530\] final_design.cpu.reg_window\[562\] net818
+ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout880_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12317__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07019_ net546 _01968_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__or2_1
X_10030_ _02837_ _04352_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07932__S net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11828__A0 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout933_X net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _06183_ net284 net405 net1698 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__a22o_1
XANTENNA__09497__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__X _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ clknet_leaf_131_clk _00951_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[708\]
+ sky130_fd_sc_hd__dfrtp_1
X_10932_ net976 _05660_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13651_ clknet_leaf_36_clk _00882_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[639\]
+ sky130_fd_sc_hd__dfrtp_1
X_10863_ _05593_ _05594_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__and2b_1
XFILLER_0_168_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12602_ net2502 net1011 net997 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1
+ vccd1 _01295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12253__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13582_ clknet_leaf_116_clk _00813_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[570\]
+ sky130_fd_sc_hd__dfrtp_1
X_10794_ net76 net1055 vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10803__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12533_ _06258_ net503 net325 net2542 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10803__B2 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12005__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12464_ net681 _06124_ _06260_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__or3_1
X_14203_ net1272 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11415_ net1950 net223 net311 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12395_ net1906 net177 net271 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14134_ clknet_leaf_77_clk final_design.vga.h_next_count\[3\] net1254 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09447__X _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11346_ _04917_ net663 vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__nand2_1
XANTENNA__12308__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07983__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14065_ clknet_leaf_46_clk _00027_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11277_ _01939_ _05947_ _05974_ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_120_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13016_ clknet_leaf_133_clk _00247_ net1166 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10228_ final_design.uart.BAUD_counter\[10\] _05104_ net811 vssd1 vssd1 vccd1 vccd1
+ _05106_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07735__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10159_ final_design.VGA_data_control.h_count\[4\] _05050_ final_design.VGA_data_control.h_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__a21oi_1
Xhold2 final_design.cpu.reg_window\[0\] vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07842__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11872__B net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12087__A3 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13918_ clknet_leaf_149_clk _01149_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[906\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12492__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10488__B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13849_ clknet_leaf_166_clk _01080_ net1105 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[837\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11047__A1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07370_ final_design.cpu.reg_window\[579\] final_design.cpu.reg_window\[611\] net942
+ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
XANTENNA__12244__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09645__D1 _04558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12195__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09040_ _03694_ _03729_ _03692_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09430__B1_N _04231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07649__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 final_design.cpu.reg_window\[238\] vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 final_design.cpu.reg_window\[747\] vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold424 final_design.cpu.reg_window\[682\] vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06921__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold435 final_design.cpu.reg_window\[475\] vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 final_design.cpu.reg_window\[47\] vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold457 final_design.uart.BAUD_counter\[16\] vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold468 final_design.cpu.reg_window\[909\] vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11539__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09942_ _03421_ _04149_ _03390_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__a21oi_1
Xhold479 final_design.cpu.reg_window\[451\] vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout904 net906 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout915 net916 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__buf_4
XANTENNA__07318__A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout926 net933 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
Xfanout937 net938 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__clkbuf_4
X_09873_ net480 _04109_ _04308_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__or3_1
Xfanout948 net956 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout294_A _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout959 net962 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _03660_ _03773_ _03661_ _03659_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__o211a_1
Xhold1102 final_design.cpu.reg_window\[54\] vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 final_design.cpu.reg_window\[34\] vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A _05167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 final_design.cpu.reg_window\[289\] vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 final_design.cpu.reg_window\[107\] vssd1 vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 final_design.cpu.reg_window\[612\] vssd1 vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09533__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08755_ _01366_ _02297_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__nor2_1
Xhold1157 final_design.cpu.reg_window\[377\] vssd1 vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 final_design.cpu.reg_window\[804\] vssd1 vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 final_design.cpu.reg_window\[801\] vssd1 vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12078__A3 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__A1 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ final_design.cpu.reg_window\[539\] final_design.cpu.reg_window\[571\] net881
+ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__mux2_1
XANTENNA__12483__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08686_ _02325_ net488 vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10398__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07637_ _02584_ _02585_ _02586_ _02587_ net694 net713 vssd1 vssd1 vccd1 vccd1 _02588_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_120_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout726_A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12235__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06892__A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ final_design.cpu.reg_window\[415\] final_design.cpu.reg_window\[447\] net841
+ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11589__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09307_ net493 _04225_ _04205_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__or3b_1
X_06519_ final_design.reqhand.instruction\[0\] final_design.reqhand.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07499_ _02032_ _02449_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__or2_1
XANTENNA__09651__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12250__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1256_X net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07199__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09238_ _04144_ _04153_ _04154_ _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_161_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09169_ _03631_ _03649_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11200_ _03995_ _05907_ net742 vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__mux2_1
XANTENNA__07927__S net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11957__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09954__A2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ _06121_ net504 _06270_ net1947 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__a22o_1
XANTENNA__08612__A _02294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11449__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ _05841_ _05844_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__nand2_2
Xhold980 final_design.cpu.reg_window\[865\] vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold991 final_design.cpu.reg_window\[584\] vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ _05783_ _05784_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__nor2_1
XANTENNA__07717__A1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ net472 _04834_ _04931_ net484 vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__o211a_1
XANTENNA__07662__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12069__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__S net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11964_ _06166_ net281 net404 net1805 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__a22o_1
XANTENNA__12474__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13703_ clknet_leaf_9_clk _00934_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[691\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10915_ _05643_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_80_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11895_ net216 net1752 net275 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output109_A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__S net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12226__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13634_ clknet_leaf_23_clk _00865_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[622\]
+ sky130_fd_sc_hd__dfrtp_1
X_10846_ net46 _05566_ _05575_ _05577_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__and4_1
XANTENNA__08493__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13565_ clknet_leaf_32_clk _00796_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[553\]
+ sky130_fd_sc_hd__dfrtp_1
X_10777_ net75 _05486_ _05512_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12241__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12516_ _06178_ net343 net327 net1556 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13496_ clknet_leaf_135_clk _00727_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[484\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12447_ net1937 net206 net335 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11201__A1 _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08602__C1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12378_ net1687 net207 net271 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__mux2_1
X_14117_ clknet_leaf_42_clk _01314_ net1153 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_11329_ _01756_ net649 _06021_ net652 _06020_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14048_ clknet_leaf_48_clk _00009_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11883__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06870_ _01485_ _01489_ _01495_ _01820_ _01502_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a41o_4
XFILLER_0_98_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07572__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11268__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ final_design.cpu.reg_window\[449\] final_design.cpu.reg_window\[481\] net849
+ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12465__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08133__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09640__X _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08471_ net612 _03415_ _03417_ net533 vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__o211a_1
XANTENNA__09881__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11822__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07422_ final_design.cpu.reg_window\[129\] final_design.cpu.reg_window\[161\] net931
+ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__mux2_1
XANTENNA__12217__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12768__A1 final_design.VGA_adr\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10946__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13006__RESET_B net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07353_ final_design.cpu.reg_window\[387\] final_design.cpu.reg_window\[419\] net943
+ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__mux2_1
XANTENNA__09094__C1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08436__A2 _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__A3 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11123__A _02095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11440__A1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07284_ final_design.cpu.reg_window\[710\] final_design.cpu.reg_window\[742\] net913
+ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09023_ _03687_ _03733_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout307_A net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 final_design.cpu.reg_window\[198\] vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_1__f_clk_X clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06651__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09936__A2 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold221 net135 vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 final_design.VGA_data_control.ready_data\[17\] vssd1 vssd1 vccd1 vccd1 net1585
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09492__S0 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold243 net133 vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold254 final_design.cpu.reg_window\[197\] vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 net162 vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold276 final_design.cpu.reg_window\[723\] vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1216_A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold287 final_design.cpu.reg_window\[227\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout701 _01753_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_4
Xfanout712 net714 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_4
Xhold298 final_design.cpu.reg_window\[855\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _03424_ _03561_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__nor2_1
Xfanout723 net724 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout734 _01493_ vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_2
XANTENNA_fanout676_A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 _01490_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_123_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 net757 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_8
Xfanout767 _01426_ vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_4
X_09856_ _04773_ _04774_ _04220_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__a21o_1
Xfanout778 net782 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_8
Xfanout789 net790 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09263__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ final_design.CPU_instr_adr\[22\] _01755_ vssd1 vssd1 vccd1 vccd1 _03758_
+ sky130_fd_sc_hd__xnor2_1
X_09787_ _03388_ _03421_ _04149_ _03389_ _03358_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__a311o_1
X_06999_ final_design.cpu.reg_window\[207\] final_design.cpu.reg_window\[239\] net907
+ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout843_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11259__A1 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ final_design.CPU_instr_adr\[11\] _02097_ vssd1 vssd1 vccd1 vccd1 _03689_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_96_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ _01999_ _02029_ _02061_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ _05400_ _05418_ _05419_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12208__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ net432 net584 _06198_ net297 net1759 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__a32o_1
XFILLER_0_83_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10631_ _05349_ _05368_ _05369_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__and3_1
XFILLER_0_166_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12223__A3 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13350_ clknet_leaf_3_clk _00581_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[338\]
+ sky130_fd_sc_hd__dfrtp_1
X_10562_ _05306_ _05308_ net1669 net1045 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12301_ net2053 net240 net366 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__mux2_1
XANTENNA__14117__Q final_design.reqhand.data_from_UART\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_134_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11982__A2 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13281_ clknet_leaf_151_clk _00512_ net1116 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[269\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10493_ net979 _05240_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09388__A0 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11320__X _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09438__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12232_ net588 _06162_ net515 net374 net2107 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_20_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11687__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11195__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08286__S1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11734__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ _06117_ _06260_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__or2_1
X_14209__1278 vssd1 vssd1 vccd1 vccd1 _14209__1278/HI net1278 sky130_fd_sc_hd__conb_1
XFILLER_0_20_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ _05065_ _05082_ _05832_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_9_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12094_ net681 _06091_ net519 vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__and3_2
XANTENNA__08038__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11907__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11045_ final_design.CPU_instr_adr\[28\] _03829_ net1072 vssd1 vssd1 vccd1 vccd1
+ _05769_ sky130_fd_sc_hd__mux2_1
XANTENNA__08488__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09173__A _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12996_ net1338 _00227_ net1159 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07549__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12__f_clk_X clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09901__A _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11947_ _06148_ net284 net409 net2404 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13170__RESET_B net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06677__A1 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ _06112_ net292 net523 net2218 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__a22o_1
XANTENNA__08517__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13617_ clknet_leaf_105_clk _00848_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[605\]
+ sky130_fd_sc_hd__dfrtp_1
X_10829_ _01385_ _05539_ _05544_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_67_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11422__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13548_ clknet_leaf_125_clk _00779_ net1196 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[536\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09091__A2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11973__A2 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13479_ clknet_leaf_9_clk _00710_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[467\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07567__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07971_ _02918_ _02919_ _02920_ _02921_ net686 net700 vssd1 vssd1 vccd1 vccd1 _02922_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_71_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11817__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ _03068_ _03101_ _04627_ net448 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_143_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06922_ _01869_ _01870_ _01871_ _01872_ net774 net795 vssd1 vssd1 vccd1 vccd1 _01873_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_143_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12061__X _06264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__A final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ net481 _04258_ _04259_ net494 vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__o31a_1
X_06853_ final_design.cpu.reg_window\[788\] final_design.cpu.reg_window\[820\] net949
+ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__mux2_1
XANTENNA__13940__RESET_B net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06500__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09572_ net474 _04260_ _04490_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10022__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06784_ final_design.cpu.reg_window\[150\] final_design.cpu.reg_window\[182\] net902
+ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__mux2_1
X_08523_ _03470_ _03471_ _03472_ _03473_ net693 net712 vssd1 vssd1 vccd1 vccd1 _03474_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08657__A2 _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__S1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout257_A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11405__X _06089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08454_ final_design.cpu.reg_window\[772\] final_design.cpu.reg_window\[804\] net860
+ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07405_ _02343_ _02344_ _02355_ net898 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_108_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08385_ final_design.cpu.reg_window\[198\] final_design.cpu.reg_window\[230\] net831
+ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__mux2_1
XANTENNA__12205__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1166_A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08146__B _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07050__B _02000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ _02283_ _02284_ _02285_ _02286_ net783 net802 vssd1 vssd1 vccd1 vccd1 _02287_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11964__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11788__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout212_X net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07267_ final_design.cpu.reg_window\[454\] final_design.cpu.reg_window\[486\] net917
+ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__mux2_1
XANTENNA__12383__S net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11140__X _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__Y _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09006_ _03791_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_115_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09258__A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07198_ final_design.cpu.reg_window\[585\] final_design.cpu.reg_window\[617\] net923
+ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_167_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11177__B1 _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout793_A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07049__Y _02000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__A3 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1121_X net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_131_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1219_X net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout960_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 net521 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_4
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout542 _02091_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_2
X_09908_ _04808_ _04826_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__xnor2_1
Xfanout553 _01784_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_4
Xfanout564 _06238_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_2
Xfanout575 net576 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_4
Xfanout586 net588 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_4
X_09839_ _04754_ _04757_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__nand2_1
Xfanout597 _05868_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08896__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout846_X net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ clknet_leaf_83_clk _00088_ net1248 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07940__S net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11801_ net2354 net413 net284 _06032_ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_140_Left_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11315__X _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11732_ net580 net422 _06224_ net296 net1784 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__a32o_1
XANTENNA__10455__A2 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11652__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08337__A _02186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10586__B final_design.VGA_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11663_ net180 net641 vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13402_ clknet_leaf_152_clk _00633_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[390\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10614_ _05357_ net970 net973 _05356_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_92_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ net183 net645 vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__and2_1
XANTENNA__07703__S0 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11955__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13333_ clknet_leaf_24_clk _00564_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[321\]
+ sky130_fd_sc_hd__dfrtp_1
X_10545_ _05290_ _05291_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_130_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07387__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13264_ clknet_leaf_115_clk _00495_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[252\]
+ sky130_fd_sc_hd__dfrtp_1
X_10476_ net976 _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__or2_1
XANTENNA__11168__A0 final_design.reqhand.data_from_UART\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08072__A _01881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ net566 _06143_ net505 net376 net1637 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__a32o_1
XFILLER_0_60_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13195_ clknet_leaf_15_clk _00426_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[183\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12146_ net222 net2243 net387 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12077_ net569 _05973_ net506 net392 net1865 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__a32o_1
XFILLER_0_60_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08336__B2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ _05731_ _05749_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08431__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06898__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09631__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire225_A _05897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12979_ clknet_leaf_68_clk _00004_ net1221 vssd1 vssd1 vccd1 vccd1 wb_manage.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11225__X _05930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08195__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12199__A2 _06127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ final_design.cpu.reg_window\[911\] final_design.cpu.reg_window\[943\] net824
+ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06990__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08534__X _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07121_ _02068_ _02069_ _02070_ _02071_ net783 net802 vssd1 vssd1 vccd1 vccd1 _02072_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11946__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_121_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07052_ final_design.cpu.reg_window\[333\] final_design.cpu.reg_window\[365\] net917
+ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XANTENNA__10017__A _03627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10382__B2 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07783__C1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12659__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07954_ _01909_ net609 vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__nand2_1
XANTENNA__11774__C net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06905_ _01850_ _01854_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__or2_1
XFILLER_0_173_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07885_ _02833_ _02835_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout374_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ _04072_ _04540_ _04541_ _04542_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__or4_1
X_06836_ final_design.data_from_mem\[21\] net983 _01786_ vssd1 vssd1 vccd1 vccd1 _01787_
+ sky130_fd_sc_hd__a21oi_2
XANTENNA__11882__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06984__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09555_ net448 _04472_ _04470_ net737 vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__o211ai_4
X_06767_ net896 _01710_ _01716_ _01703_ _01704_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__a32o_2
XANTENNA__09288__C1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12378__S net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A _06157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ net625 _03450_ _03451_ _02326_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__a211o_1
XANTENNA__11634__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ _01566_ net455 _04207_ net468 vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__a211o_1
XFILLER_0_148_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06698_ _01645_ _01646_ _01647_ _01648_ net785 net803 vssd1 vssd1 vccd1 vccd1 _01649_
+ sky130_fd_sc_hd__mux4_1
X_14208__1277 vssd1 vssd1 vccd1 vccd1 _14208__1277/HI net1277 sky130_fd_sc_hd__conb_1
XFILLER_0_148_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08437_ net534 _03386_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout806_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08368_ _03315_ _03316_ _03317_ _03318_ net686 net702 vssd1 vssd1 vccd1 vccd1 _03319_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11398__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07319_ _02268_ _02269_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__and2b_1
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_112_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08299_ net726 _03249_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__nor2_1
XANTENNA__11311__A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10330_ net1516 net1025 net1002 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1
+ vccd1 _00087_ sky130_fd_sc_hd__a22o_1
XANTENNA__07161__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10261_ net1728 _05124_ _05126_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06899__X _01850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ _06202_ net282 net400 net2353 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__a22o_1
XANTENNA__12362__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13862__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ final_design.uart.BAUD_counter\[2\] final_design.uart.BAUD_counter\[7\] final_design.uart.BAUD_counter\[6\]
+ final_design.uart.BAUD_counter\[3\] vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__or4b_1
XANTENNA__08620__A _02127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__B2 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11457__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout350 net351 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_4
Xfanout361 net363 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_6
XANTENNA__09515__A0 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07236__A _02185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout372 net373 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11322__A0 _04597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13951_ clknet_leaf_135_clk _01182_ net1167 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[939\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout383 _06269_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_4
Xfanout394 net395 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_8
X_12902_ clknet_leaf_68_clk _00140_ net1221 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__dfrtp_1
X_13882_ clknet_leaf_163_clk _01113_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[870\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11873__B2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12833_ net1394 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10428__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12764_ _05039_ _06382_ _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11715_ net195 net634 vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12695_ final_design.VGA_data_control.v_count\[5\] _06335_ vssd1 vssd1 vccd1 vccd1
+ _06336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11920__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input92_X net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11646_ net435 net587 _06180_ net301 net1600 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_42_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11928__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 mem_adr_start[0] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
XFILLER_0_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11577_ net569 net421 _06144_ net303 net2028 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_103_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
Xinput47 mem_adr_start[1] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_1
XFILLER_0_13_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput58 mem_adr_start[2] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_1
XANTENNA__06804__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11221__A _04744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13316_ clknet_leaf_100_clk _00547_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[304\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput69 memory_size[10] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_4
X_10528_ final_design.CPU_instr_adr\[4\] _05275_ net1068 vssd1 vssd1 vccd1 vccd1 _05276_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold809 final_design.cpu.reg_window\[961\] vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13247_ clknet_leaf_134_clk _00478_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[235\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10459_ net1445 net1048 _05213_ net248 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07845__S net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12353__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ clknet_leaf_164_clk _00409_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[166\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11875__B net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10364__B2 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _05840_ _05841_ _05858_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__and3_2
XANTENNA__08309__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07670_ _02617_ _02618_ _02619_ _02620_ net687 net708 vssd1 vssd1 vccd1 vccd1 _02621_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_88_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11864__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07580__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06966__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ final_design.cpu.reg_window\[347\] final_design.cpu.reg_window\[379\] net961
+ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09340_ _04078_ _04102_ net469 vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__a21oi_1
X_06552_ _01484_ _01488_ net747 _01494_ _01501_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__o41a_1
XANTENNA__11616__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09271_ net80 net81 _04189_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__or3_2
XFILLER_0_59_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06483_ final_design.cpu.reg_window\[158\] final_design.cpu.reg_window\[190\] net928
+ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11830__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08222_ _03169_ _03170_ _03171_ _03172_ net691 net711 vssd1 vssd1 vccd1 vccd1 _03173_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_114_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07391__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06924__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07048__A1 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11919__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12041__A1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08153_ _01968_ net617 vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_151_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07104_ final_design.cpu.reg_window\[524\] final_design.cpu.reg_window\[556\] net928
+ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08084_ _02803_ _03034_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07035_ final_design.cpu.reg_window\[910\] final_design.cpu.reg_window\[942\] net925
+ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10970__A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12344__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__B2 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__A1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08986_ _03745_ _03746_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07937_ final_design.cpu.reg_window\[726\] final_design.cpu.reg_window\[758\] net819
+ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07868_ final_design.cpu.reg_window\[788\] final_design.cpu.reg_window\[820\] net876
+ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
XANTENNA__08586__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08181__C1 _01966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09607_ net264 _04516_ _04522_ _04525_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__and4_1
X_06819_ _01766_ _01767_ _01768_ _01769_ net789 net806 vssd1 vssd1 vccd1 vccd1 _01770_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_27_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07799_ net729 _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout923_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08159__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09538_ net552 net551 net549 net548 net453 net462 vssd1 vssd1 vccd1 vccd1 _04457_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_167_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09469_ _04385_ _04387_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12280__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11740__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ _05840_ _05842_ _06117_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__nor3_1
XFILLER_0_136_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12480_ _06140_ net345 net331 net2369 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11431_ net1944 _06017_ net313 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14150_ clknet_leaf_80_clk _01324_ net1249 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11362_ net664 _06048_ _06050_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__or3_1
XFILLER_0_105_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06798__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13101_ clknet_leaf_104_clk _00332_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11791__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10313_ final_design.VGA_data_control.state\[0\] _01394_ final_design.VGA_data_control.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14081_ clknet_leaf_71_clk _01278_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11293_ net426 net571 _05990_ net315 net1998 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13032_ clknet_leaf_125_clk _00263_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12335__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input52_A mem_adr_start[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ final_design.uart.BAUD_counter\[16\] _05114_ net809 vssd1 vssd1 vccd1 vccd1
+ _05116_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11695__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10346__B2 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1103 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__clkbuf_2
Xfanout1112 net1118 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_4
X_10175_ final_design.uart.bits_received\[1\] final_design.uart.bits_received\[2\]
+ _05064_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__nor3_1
Xfanout1123 net1124 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__clkbuf_4
Xfanout1134 net1137 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__buf_2
XFILLER_0_100_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1145 net1156 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12099__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1156 net1164 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__clkbuf_4
Xfanout1167 net1168 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__buf_2
Xfanout180 _06074_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
Xfanout1178 net1181 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1189 net100 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkbuf_4
Xfanout191 _06038_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
X_13934_ clknet_leaf_119_clk _01165_ net1199 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[922\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12996__RESET_B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08496__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13865_ clknet_leaf_87_clk _01096_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[853\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12816_ net1365 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_83_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13796_ clknet_leaf_106_clk _01027_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[784\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12747_ final_design.VGA_adr\[4\] net808 vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12678_ _06326_ net1497 net993 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11629_ net211 net639 vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08322__S0 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13784__RESET_B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10585__A1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold606 final_design.cpu.reg_window\[342\] vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 final_design.cpu.reg_window\[848\] vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11782__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold628 final_design.cpu.reg_window\[843\] vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold639 final_design.cpu.reg_window\[664\] vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_59_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10337__B2 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14207__1276 vssd1 vssd1 vccd1 vccd1 _14207__1276/HI net1276 sky130_fd_sc_hd__conb_1
X_08840_ final_design.CPU_instr_adr\[14\] _03790_ vssd1 vssd1 vccd1 vccd1 _03791_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_85_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08771_ _03704_ _03721_ _03703_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06986__Y _01937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11825__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ _02670_ _02671_ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__or2_2
XANTENNA__06919__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10949__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08702__A1 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07653_ net613 _02602_ _02577_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06604_ final_design.cpu.reg_window\[796\] final_design.cpu.reg_window\[828\] net954
+ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07584_ final_design.cpu.reg_window\[799\] final_design.cpu.reg_window\[831\] net841
+ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09323_ _04241_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__inv_2
X_06535_ _01456_ _01465_ _01474_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__nor3_1
XFILLER_0_164_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12262__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout337_A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ _02574_ _02606_ _04171_ _02641_ _02575_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__a311o_1
XANTENNA_fanout1079_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06466_ final_design.reqhand.instruction\[17\] net984 vssd1 vssd1 vccd1 vccd1 _01417_
+ sky130_fd_sc_hd__or2_1
XANTENNA__06654__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12953__Q net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ final_design.cpu.reg_window\[590\] final_design.cpu.reg_window\[622\] net853
+ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11132__Y _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09185_ _04102_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout504_A _06264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1246_A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08136_ final_design.cpu.reg_window\[717\] final_design.cpu.reg_window\[749\] net832
+ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__mux2_1
XANTENNA__10576__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10576__B2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07441__A1 final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11796__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ final_design.cpu.reg_window\[594\] final_design.cpu.reg_window\[626\] net818
+ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12391__S net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07018_ _01966_ _01968_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10328__B2 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ net630 _03906_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11980_ _06182_ net278 net404 net2013 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__a22o_1
X_10931_ net972 _05656_ _05659_ net968 vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10862_ _05569_ _05586_ _05587_ _05592_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__or4_1
X_13650_ clknet_leaf_44_clk _00881_ net1150 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[638\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12601_ net2413 net1010 net996 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1
+ vccd1 _01294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13581_ clknet_leaf_139_clk _00812_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[569\]
+ sky130_fd_sc_hd__dfrtp_1
X_10793_ net76 net1055 vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__and2_1
XANTENNA__11470__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12532_ _06195_ net350 net324 net2199 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12463_ net1684 net177 net336 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__mux2_1
XANTENNA__08304__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14202_ net1271 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
X_11414_ net2330 net239 net313 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__mux2_1
XANTENNA__12556__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12394_ net1685 net179 net271 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14133_ clknet_leaf_77_clk final_design.vga.h_next_count\[2\] net1254 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11345_ _01691_ net650 _06035_ net652 net663 vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07395__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07983__A2 _02929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14064_ clknet_leaf_46_clk _00026_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11276_ net743 _03927_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10319__B2 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13015_ clknet_leaf_144_clk _00246_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10227_ _05104_ _05105_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ final_design.VGA_data_control.h_count\[4\] final_design.VGA_data_control.h_count\[5\]
+ _05050_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_131_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 final_design.cpu.reg_window\[9\] vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ final_design.vga.v_current_state\[1\] final_design.vga.v_current_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_85_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07424__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13917_ clknet_leaf_13_clk _01148_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[905\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_146_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13848_ clknet_leaf_129_clk _01079_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[836\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12244__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09645__C1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13779_ clknet_leaf_34_clk _01010_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[767\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08255__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12547__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11755__A0 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 final_design.cpu.reg_window\[90\] vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold414 final_design.cpu.reg_window\[56\] vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 final_design.cpu.reg_window\[833\] vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold436 final_design.cpu.reg_window\[248\] vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold447 final_design.cpu.reg_window\[763\] vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 final_design.cpu.reg_window\[88\] vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 final_design.cpu.reg_window\[971\] vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _04719_ _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_129_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10616__A1_N net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout905 net906 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
Xfanout916 net917 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_4
Xfanout927 net929 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _03522_ _04087_ _04094_ _03520_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a221o_1
Xfanout938 net945 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_4
Xfanout949 net950 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _03660_ _03773_ _03661_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__o21a_1
Xhold1103 final_design.cpu.reg_window\[121\] vssd1 vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 final_design.cpu.reg_window\[610\] vssd1 vssd1 vccd1 vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1125 final_design.cpu.reg_window\[738\] vssd1 vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout287_A _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1136 final_design.cpu.reg_window\[99\] vssd1 vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ _03703_ _03704_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__nand2b_1
Xhold1147 final_design.cpu.reg_window\[295\] vssd1 vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 final_design.cpu.reg_window\[926\] vssd1 vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 final_design.cpu.reg_window\[908\] vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ final_design.cpu.reg_window\[603\] final_design.cpu.reg_window\[635\] net881
+ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__mux2_1
XANTENNA__12948__Q net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08685_ _03486_ _03487_ _03520_ _03521_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__o22a_1
XFILLER_0_136_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout454_A net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1196_A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07636_ final_design.cpu.reg_window\[156\] final_design.cpu.reg_window\[188\] net874
+ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12235__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12386__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07567_ final_design.cpu.reg_window\[479\] final_design.cpu.reg_window\[511\] net845
+ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout621_A _02513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout242_X net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09306_ net474 net465 net530 vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11143__X _05858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06518_ _01466_ _01467_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07498_ _02067_ _02101_ _02446_ _02065_ _02033_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__o311a_1
XANTENNA__08165__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09237_ _04141_ _04155_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__or2_1
X_06449_ final_design.VGA_data_control.v_count\[7\] final_design.VGA_data_control.v_count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__nand2_1
X_12801__32 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__inv_2
XFILLER_0_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12538__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09168_ _03631_ net666 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__nor2_4
XFILLER_0_146_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11746__A0 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08119_ _03067_ _03069_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09099_ final_design.CPU_instr_adr\[3\] net1031 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__xor2_1
XFILLER_0_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11957__C net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08612__B net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11130_ _05842_ _05843_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__nor2_2
XFILLER_0_31_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold970 final_design.cpu.reg_window\[535\] vssd1 vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold981 final_design.cpu.reg_window\[277\] vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ _05763_ _05765_ _05779_ _05782_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__o211a_1
Xhold992 final_design.cpu.reg_window\[831\] vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
X_10012_ net475 _04930_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__nand2_1
XANTENNA__08914__B2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11465__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ _06165_ net279 net404 net1603 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_83_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13702_ clknet_leaf_170_clk _00933_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[690\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ net50 _05642_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11894_ net218 net2120 net274 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10845_ _05566_ _05575_ _05577_ net46 vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__a31oi_2
X_13633_ clknet_leaf_157_clk _00864_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[621\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12226__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14206__1275 vssd1 vssd1 vccd1 vccd1 _14206__1275/HI net1275 sky130_fd_sc_hd__conb_1
XFILLER_0_55_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10776_ _05510_ _05511_ _05486_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_137_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13564_ clknet_leaf_151_clk _00795_ net1116 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[552\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11985__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09642__A2 _04559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12515_ _06177_ net346 net327 net1862 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__a22o_1
X_13495_ clknet_leaf_143_clk _00726_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[483\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12529__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12446_ net1814 net207 net336 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11201__A2 _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12377_ net1592 net210 net270 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__mux2_1
XANTENNA__07405__B2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08602__B1 _03524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14116_ clknet_leaf_52_clk net1415 net1151 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11328_ final_design.data_from_mem\[22\] net236 net234 vssd1 vssd1 vccd1 vccd1 _06021_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__10960__A1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10960__B2 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14047_ clknet_leaf_48_clk _00008_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11259_ final_design.data_from_mem\[14\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1
+ _05960_ sky130_fd_sc_hd__a21o_2
XFILLER_0_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09193__X _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12940__RESET_B net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12331__Y _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12060__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08118__C1 _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12465__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_74_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_35_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08470_ _02294_ net496 vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__or2_2
XFILLER_0_148_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07421_ final_design.cpu.reg_window\[193\] final_design.cpu.reg_window\[225\] net931
+ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08516__S0 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12768__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07352_ final_design.cpu.reg_window\[451\] final_design.cpu.reg_window\[483\] net943
+ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11976__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07283_ final_design.cpu.reg_window\[518\] final_design.cpu.reg_window\[550\] net913
+ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09022_ _02067_ _02447_ _03953_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11728__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold200 final_design.cpu.reg_window\[711\] vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold211 final_design.cpu.reg_window\[467\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold222 final_design.cpu.reg_window\[860\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold233 final_design.VGA_data_control.ready_data\[8\] vssd1 vssd1 vccd1 vccd1 net1586
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09492__S1 _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold244 final_design.cpu.reg_window\[237\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold255 final_design.cpu.reg_window\[800\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold266 final_design.reqhand.instruction\[0\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 final_design.cpu.reg_window\[229\] vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold288 final_design.cpu.reg_window\[575\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 final_design.cpu.reg_window\[557\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout702 net703 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__clkbuf_8
X_09924_ net264 _04837_ _04841_ _04842_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__and4_1
Xfanout713 net714 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout724 _01721_ vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1111_A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout735 _01493_ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07763__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1209_A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout746 net748 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_2
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout757 _01438_ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_8
X_09855_ net603 _04266_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__nand2_1
XANTENNA__11900__A0 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 _01426_ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__buf_2
XANTENNA_fanout571_A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout779 net780 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08806_ _03754_ _03756_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__nor2_1
X_06998_ final_design.cpu.reg_window\[15\] final_design.cpu.reg_window\[47\] net907
+ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__mux2_1
X_09786_ _03391_ _04149_ _04150_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__o21ai_1
X_08737_ final_design.CPU_instr_adr\[11\] _02097_ vssd1 vssd1 vccd1 vccd1 _03688_
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_65_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout836_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08668_ _01463_ _01484_ _03618_ _01486_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09872__A2 _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12208__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07619_ net893 _02569_ _02558_ _02557_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__o2bb2a_2
X_08599_ net891 _03542_ _03548_ _03535_ _03536_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__a32o_4
XFILLER_0_113_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10630_ _05368_ _05369_ _05349_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09085__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11967__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10561_ net1018 _05304_ _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__or3_1
XANTENNA__08832__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12300_ net2214 net227 net366 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07938__S net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13280_ clknet_leaf_35_clk _00511_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[268\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10492_ net978 _05241_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08623__A _02185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12231_ _06161_ net501 net373 net2436 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_20_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09388__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09438__B _04190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11195__A1 _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12162_ _06117_ _06260_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__nor2_1
X_11113_ final_design.uart.bits_received\[0\] final_design.uart.bits_received\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_9_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12093_ net580 _06090_ net511 net393 net1641 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__a32o_1
XANTENNA__12144__A0 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07673__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ final_design.CPU_instr_adr\[28\] net1014 _05767_ net1054 net975 vssd1 vssd1
+ vccd1 vccd1 _05768_ sky130_fd_sc_hd__o221a_1
XANTENNA__08899__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__A1 _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09173__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12447__A1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12995_ net1337 _00226_ net1159 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07549__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11946_ _06147_ net278 net408 net2046 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11877_ _06111_ net291 net522 net1854 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__a22o_1
X_13616_ clknet_leaf_104_clk _00847_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[604\]
+ sky130_fd_sc_hd__dfrtp_1
X_10828_ _05559_ _05561_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08009__S net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13547_ clknet_leaf_16_clk _00778_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[535\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10759_ _05483_ _05493_ _05495_ net42 vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13478_ clknet_leaf_171_clk _00709_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[466\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12792__23 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__inv_2
X_12429_ final_design.cpu.reg_window\[895\] net340 vssd1 vssd1 vccd1 vccd1 _06281_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07970_ final_design.cpu.reg_window\[785\] final_design.cpu.reg_window\[817\] net836
+ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08339__C1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07583__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06921_ final_design.cpu.reg_window\[914\] final_design.cpu.reg_window\[946\] net901
+ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_0__f_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_06852_ final_design.cpu.reg_window\[852\] final_design.cpu.reg_window\[884\] net949
+ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__mux2_1
X_09640_ _04486_ _04489_ net480 vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_160_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09571_ net475 _04489_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__nand2_1
XANTENNA__12438__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06783_ final_design.cpu.reg_window\[214\] final_design.cpu.reg_window\[246\] net902
+ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__mux2_1
XANTENNA__10022__B _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk
+ sky130_fd_sc_hd__clkbuf_8
X_08522_ final_design.cpu.reg_window\[898\] final_design.cpu.reg_window\[930\] net865
+ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__mux2_1
XANTENNA__11833__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13980__RESET_B net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08453_ final_design.cpu.reg_window\[836\] final_design.cpu.reg_window\[868\] net859
+ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__mux2_1
XANTENNA__09530__C _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07404_ _02349_ _02354_ net762 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08384_ final_design.cpu.reg_window\[6\] final_design.cpu.reg_window\[38\] net831
+ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11949__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07335_ final_design.cpu.reg_window\[900\] final_design.cpu.reg_window\[932\] net940
+ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10973__A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout417_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1159_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07266_ final_design.cpu.reg_window\[262\] final_design.cpu.reg_window\[294\] net914
+ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__mux2_1
XANTENNA__11788__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09005_ final_design.CPU_instr_adr\[14\] _03790_ vssd1 vssd1 vccd1 vccd1 _03939_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07197_ net760 _02147_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__or2_1
XANTENNA__11177__A1 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout786_A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14086__RESET_B net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08589__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout510 net513 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09274__A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07346__X _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout521 net523 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_4
Xfanout532 _02356_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__clkbuf_4
X_09907_ _04072_ _04824_ _04810_ net738 vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__o211a_1
Xfanout543 _02058_ vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_2
X_14205__1274 vssd1 vssd1 vccd1 vccd1 _14205__1274/HI net1274 sky130_fd_sc_hd__conb_1
XANTENNA__12677__B2 final_design.data_from_mem\[26\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout953_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout554 _01750_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 _05869_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_8
Xfanout576 _05868_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_2
Xfanout587 net588 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_2
X_09838_ net493 _04435_ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a21o_1
Xfanout598 net600 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ _03588_ net442 net439 _03587_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_38_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11743__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11800_ net2533 net412 _06236_ net425 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__a22o_1
XANTENNA__09721__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11731_ net178 net635 vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__and2_1
XANTENNA__11652__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08337__B net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11662_ net436 net590 _06188_ net301 net1584 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_25_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13401_ clknet_leaf_165_clk _00632_ net1085 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[389\]
+ sky130_fd_sc_hd__dfrtp_1
X_10613_ final_design.CPU_instr_adr\[8\] _03988_ net1071 vssd1 vssd1 vccd1 vccd1 _05357_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11593_ net596 net424 _06152_ net306 net1536 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__a32o_1
XFILLER_0_153_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12601__B2 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11331__X _06024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07668__S net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input82_A memory_size[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10544_ net94 final_design.VGA_adr\[2\] _05289_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__and3_1
X_13332_ clknet_leaf_103_clk _00563_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[320\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07703__S1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12871__Q final_design.data_from_mem\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10475_ net79 net971 net969 final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1
+ _05226_ sky130_fd_sc_hd__o22a_1
XFILLER_0_161_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13263_ clknet_leaf_92_clk _00494_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[251\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09168__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__A1 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08072__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08569__C1 _02390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12214_ net571 _06142_ net507 net376 net2147 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__a32o_1
XANTENNA__11210__C _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13194_ clknet_leaf_1_clk _00425_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[182\]
+ sky130_fd_sc_hd__dfrtp_1
X_12145_ net205 net2424 net384 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12076_ net2548 net393 net500 _05966_ vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__a22o_1
X_11027_ net1016 _05750_ _05751_ net1046 net1379 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__a32o_1
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10123__A final_design.VGA_data_control.v_count\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_155_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13738__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09190__Y _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10410__X _05188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12978_ clknet_leaf_69_clk _00003_ net1221 vssd1 vssd1 vccd1 vccd1 wb_manage.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_47_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08195__S1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11929_ _06131_ net279 net408 net2282 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10851__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12199__A3 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06990__B _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07120_ final_design.cpu.reg_window\[395\] final_design.cpu.reg_window\[427\] net938
+ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07578__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07051_ _01996_ _02000_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12356__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10017__B _03649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XANTENNA__11828__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06586__A1 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06511__A final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ _01910_ net617 vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__nor2_1
XANTENNA__12659__B2 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06904_ _01850_ _01854_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__and2_1
X_07884_ net608 _02830_ _02805_ _01815_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__o211a_1
XANTENNA__11331__A1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ _04536_ _04537_ _04538_ _04534_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__a31o_1
X_06835_ final_design.reqhand.instruction\[21\] net982 vssd1 vssd1 vccd1 vccd1 _01786_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11882__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_A _06275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09554_ net448 _04472_ _04470_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__o21ai_1
X_06766_ net896 _01710_ _01716_ _01703_ _01704_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__a32oi_4
XANTENNA__06657__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09288__B1 _03524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11095__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ net614 _03450_ _03452_ _02326_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__o211ai_1
X_06697_ final_design.cpu.reg_window\[921\] final_design.cpu.reg_window\[953\] net941
+ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__mux2_1
X_09485_ net530 net459 _04203_ net464 vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__a211o_1
XANTENNA__11634__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout534_A net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08436_ net621 _03384_ _03385_ net534 vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_19_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11799__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12394__S net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08367_ final_design.cpu.reg_window\[519\] final_design.cpu.reg_window\[551\] net856
+ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout701_A _01753_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11398__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07318_ net535 _02267_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08298_ _03245_ _03246_ _03247_ _03248_ net688 net709 vssd1 vssd1 vccd1 vccd1 _03249_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07697__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11311__B _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07249_ final_design.cpu.reg_window\[839\] final_design.cpu.reg_window\[871\] net937
+ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12347__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ final_design.uart.BAUD_counter\[22\] _05124_ net809 vssd1 vssd1 vccd1 vccd1
+ _05126_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07449__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11738__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ net1065 _01392_ _05080_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 net342 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_4
Xfanout351 net352 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09515__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout362 net363 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_8
Xfanout373 net375 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07236__B _02186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13950_ clknet_leaf_149_clk _01181_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[938\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout384 net385 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_8
Xfanout395 _06263_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_4
X_12901_ clknet_leaf_68_clk _00139_ net1221 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dfrtp_1
X_13881_ clknet_leaf_161_clk _01112_ net1085 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[869\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11873__A2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11473__S net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12832_ net1363 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12866__Q final_design.data_from_mem\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12763_ _06339_ _06392_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10833__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11714_ net438 net595 _06215_ net298 net1833 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12694_ _01369_ final_design.VGA_data_control.v_count\[6\] _06334_ vssd1 vssd1 vccd1
+ vccd1 _06335_ sky130_fd_sc_hd__a21o_1
XANTENNA__10884__Y _05615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06501__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11645_ net198 net640 vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_42_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09179__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input85_X net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08083__A _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11576_ net200 net642 vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__and2_1
Xinput37 mem_adr_start[10] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput48 mem_adr_start[20] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10061__A1 _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput59 mem_adr_start[30] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__buf_1
XANTENNA__11221__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13315_ clknet_leaf_5_clk _00546_ net1096 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[303\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10527_ _05273_ _05274_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12338__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09466__X _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13246_ clknet_leaf_19_clk _00477_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[234\]
+ sky130_fd_sc_hd__dfrtp_1
X_10458_ _02570_ net602 vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11010__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10389_ net813 net1016 _05175_ net1046 net1511 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__a32o_1
X_13177_ clknet_leaf_168_clk _00408_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[165\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10364__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12128_ final_design.cpu.reg_window\[608\] net386 vssd1 vssd1 vccd1 vccd1 _06267_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_165_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08309__A2 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ _05840_ _05841_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__nand2_2
XANTENNA__12510__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07612__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13572__RESET_B net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06620_ _01567_ _01570_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_172_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11077__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06551_ final_design.data_from_mem\[31\] net981 _01500_ vssd1 vssd1 vccd1 vccd1 _01502_
+ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_66_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11616__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09270_ net78 _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_103_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06482_ final_design.cpu.reg_window\[222\] final_design.cpu.reg_window\[254\] net928
+ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08221_ final_design.cpu.reg_window\[395\] final_design.cpu.reg_window\[427\] net857
+ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14204__1273 vssd1 vssd1 vccd1 vccd1 _14204__1273/HI net1273 sky130_fd_sc_hd__conb_1
XFILLER_0_145_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08152_ _03067_ _03069_ _03099_ _03100_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__o22a_1
XANTENNA__08245__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09442__B1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06506__A final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07103_ final_design.cpu.reg_window\[588\] final_design.cpu.reg_window\[620\] net928
+ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08083_ _01815_ _02832_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_9_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07034_ final_design.cpu.reg_window\[974\] final_design.cpu.reg_window\[1006\] net926
+ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__mux2_1
XANTENNA__06940__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08721__A final_design.CPU_instr_adr\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11001__B1 _05239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10355__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1024_A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ _01942_ _02455_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout484_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ net717 _02886_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07771__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12501__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout651_A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12389__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ final_design.cpu.reg_window\[852\] final_design.cpu.reg_window\[884\] net868
+ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11855__A2 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07343__Y _02294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ _04222_ _04524_ _04218_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06818_ final_design.cpu.reg_window\[405\] final_design.cpu.reg_window\[437\] net963
+ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07798_ _02745_ _02746_ _02747_ _02748_ net694 net713 vssd1 vssd1 vccd1 vccd1 _02749_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_27_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08159__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ _03585_ _03589_ _02935_ _02963_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_167_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06749_ final_design.cpu.reg_window\[215\] final_design.cpu.reg_window\[247\] net925
+ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout916_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09468_ _04193_ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08419_ _03366_ _03367_ _03368_ _03369_ net682 net704 vssd1 vssd1 vccd1 vccd1 _03370_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09399_ _02574_ net440 _04314_ _04317_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ net1949 net197 net313 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06416__A net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10043__A1 _04571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11361_ _01630_ net650 _06049_ net653 vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__a22o_1
XANTENNA__06798__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10312_ net1054 _01395_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__or2_1
X_13100_ clknet_leaf_122_clk _00331_ net1197 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14080_ clknet_leaf_71_clk _01277_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11292_ net654 net203 vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__and2_1
X_10243_ _05114_ _05115_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__nor2_1
X_13031_ clknet_leaf_8_clk _00262_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08095__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10346__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A mem_adr_start[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ final_design.uart.bits_received\[0\] final_design.uart.bits_received\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__nand2_1
Xfanout1102 net1103 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_4
Xfanout1113 net1118 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__clkbuf_2
Xfanout1124 net1128 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__clkbuf_4
Xfanout1135 net1137 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__clkbuf_4
Xfanout1146 net1149 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__clkbuf_4
Xfanout1157 net1164 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10879__Y _05610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1168 net1173 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1179 net1181 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__clkbuf_2
Xfanout181 _06074_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_2
Xfanout192 net193 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_2
X_13933_ clknet_leaf_127_clk _01164_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[921\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12299__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11846__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13864_ clknet_leaf_119_clk _01095_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[852\]
+ sky130_fd_sc_hd__dfrtp_1
X_12815_ net1380 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__clkbuf_1
X_13795_ clknet_leaf_5_clk _01026_ net1096 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[783\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _05058_ _06359_ _06366_ _06376_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__nor4_1
XFILLER_0_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07290__A_N _02239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07710__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ final_design.VGA_data_control.ready_data\[26\] net1034 net989 final_design.data_from_mem\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_13_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12559__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ net432 net583 _06171_ net301 net1745 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__a32o_1
XANTENNA__12023__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08322__S1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11231__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire560 _01596_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11559_ net430 net582 _06135_ net304 net1715 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__a32o_1
XFILLER_0_123_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold607 final_design.cpu.reg_window\[436\] vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold618 final_design.cpu.reg_window\[150\] vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07856__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold629 final_design.cpu.reg_window\[502\] vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13229_ clknet_leaf_139_clk _00460_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[217\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10337__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11534__A1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _03708_ _03720_ _03706_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07721_ _02670_ _02671_ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__nor2_1
XANTENNA__09360__C1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07652_ _01570_ net626 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__nor2_1
XANTENNA__07016__B1_N _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06603_ final_design.cpu.reg_window\[860\] final_design.cpu.reg_window\[892\] net954
+ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07583_ final_design.cpu.reg_window\[863\] final_design.cpu.reg_window\[895\] net844
+ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11841__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06534_ _01474_ _01481_ _01482_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_122_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09322_ net480 _04240_ _04236_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_122_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09663__B1 _04231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06465_ net1051 net1008 net1005 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__or3_1
X_09253_ _02574_ _02606_ _04171_ _02575_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout232_A _05858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08204_ final_design.cpu.reg_window\[654\] final_design.cpu.reg_window\[686\] net844
+ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09184_ net622 _03550_ _01536_ _02423_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__a211o_1
XFILLER_0_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12014__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08135_ final_design.cpu.reg_window\[525\] final_design.cpu.reg_window\[557\] net832
+ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12672__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1141_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11773__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1239_A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08066_ final_design.cpu.reg_window\[658\] final_design.cpu.reg_window\[690\] net818
+ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__mux2_1
XANTENNA__11796__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07619__X _02570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06670__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08451__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07017_ _01967_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout699_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1027_X net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout866_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13423__RESET_B net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ _03675_ _03750_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__xnor2_1
X_07919_ final_design.cpu.reg_window\[342\] final_design.cpu.reg_window\[374\] net822
+ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08899_ net259 _03844_ net1029 vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10930_ final_design.CPU_instr_adr\[23\] _03870_ net1071 vssd1 vssd1 vccd1 vccd1
+ _05659_ sky130_fd_sc_hd__mux2_1
XANTENNA__07006__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10861_ _05569_ _05586_ _05587_ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__o31a_1
XANTENNA__11751__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ net1405 net1010 net996 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1
+ vccd1 _01293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ clknet_leaf_125_clk _00811_ net1196 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[568\]
+ sky130_fd_sc_hd__dfrtp_1
X_10792_ _04474_ net251 vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11461__A0 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12531_ net680 net637 _06268_ net326 net1991 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08209__A1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12462_ net2511 net179 net336 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__mux2_1
XANTENNA__12005__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14201_ net1270 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_0_152_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11413_ net2403 net226 net313 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__mux2_1
XANTENNA__08304__S1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11213__B1 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12393_ net1688 net181 net273 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14132_ clknet_leaf_77_clk final_design.vga.h_next_count\[1\] net1254 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[1\] sky130_fd_sc_hd__dfrtp_2
X_11344_ final_design.data_from_mem\[24\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06035_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14063_ clknet_leaf_43_clk _00025_ net1149 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11275_ net667 _03923_ net739 vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_37_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13014_ clknet_leaf_130_clk _00245_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input48_X net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10226_ final_design.uart.BAUD_counter\[9\] _05103_ net811 vssd1 vssd1 vccd1 vccd1
+ _05105_ sky130_fd_sc_hd__o21ai_1
XANTENNA_output151_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ net1061 _05050_ _05053_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__13164__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 final_design.cpu.reg_window\[25\] vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__dlygate4sd3_1
X_14203__1272 vssd1 vssd1 vccd1 vccd1 _14203__1272/HI net1272 sky130_fd_sc_hd__conb_1
XANTENNA__09192__A _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10088_ _04997_ _05003_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_85_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11227__A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13916_ clknet_leaf_153_clk _01147_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[904\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08696__A1 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12492__A2 _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13847_ clknet_leaf_143_clk _01078_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[835\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13778_ clknet_leaf_39_clk _01009_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[766\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12729_ _06364_ _06369_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__nor2_1
XFILLER_0_167_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07656__C1 _01566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11204__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07586__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07439__X _02390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold404 final_design.cpu.reg_window\[45\] vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09367__A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold415 final_design.cpu.reg_window\[794\] vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold426 final_design.cpu.reg_window\[134\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 final_design.cpu.reg_window\[852\] vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold448 final_design.cpu.reg_window\[74\] vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold459 final_design.cpu.reg_window\[776\] vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ _03391_ _03563_ _04718_ _04046_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__o31a_1
XFILLER_0_110_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout906 net912 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_2
Xfanout917 net922 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__clkbuf_4
X_09871_ _03521_ net444 vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__nor2_1
Xfanout928 net929 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__clkbuf_4
Xfanout939 net941 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11836__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ _03663_ _03772_ _03662_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_146_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 final_design.cpu.reg_window\[119\] vssd1 vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 final_design.cpu.reg_window\[271\] vssd1 vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 final_design.cpu.reg_window\[116\] vssd1 vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 final_design.cpu.reg_window\[416\] vssd1 vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ net675 _01659_ final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1 vccd1 _03704_
+ sky130_fd_sc_hd__a21o_1
Xhold1148 final_design.cpu.reg_window\[618\] vssd1 vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout182_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1159 final_design.cpu.reg_window\[125\] vssd1 vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_124_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07704_ net729 _02654_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08684_ _03617_ net603 vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__nand2b_2
XANTENNA__12483__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07635_ final_design.cpu.reg_window\[220\] final_design.cpu.reg_window\[252\] net874
+ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10684__A_N net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1091_A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1189_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06665__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07566_ final_design.cpu.reg_window\[287\] final_design.cpu.reg_window\[319\] net845
+ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09305_ _02503_ net481 vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__nand2_1
X_06517_ _01466_ _01467_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__or2_4
XFILLER_0_1_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07497_ _02067_ _02447_ _02065_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout614_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11994__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ _03261_ _03291_ _03259_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06448_ _01397_ _01400_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09167_ _04054_ net320 vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__nand2_2
XFILLER_0_161_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08298__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_X net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11600__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09277__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08118_ net606 _03065_ _03041_ _02058_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ _02432_ _04019_ _04020_ net628 vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ final_design.cpu.reg_window\[402\] final_design.cpu.reg_window\[434\] net819
+ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13604__RESET_B net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold960 final_design.cpu.reg_window\[486\] vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold971 final_design.cpu.reg_window\[118\] vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ _05779_ _05782_ _05763_ _05765_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__a211oi_1
Xhold982 final_design.cpu.reg_window\[616\] vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 final_design.cpu.reg_window\[264\] vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ net464 _03641_ _04237_ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__a31o_1
XANTENNA__11746__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08375__B1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11962_ _06164_ net288 net406 net2176 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__a22o_1
XANTENNA__08222__S0 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__A0 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12474__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13701_ clknet_leaf_4_clk _00932_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[689\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10913_ net50 _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__and2_1
XFILLER_0_169_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11682__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11893_ net220 net2210 net275 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__mux2_1
XANTENNA__11481__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13632_ clknet_leaf_45_clk _00863_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[620\]
+ sky130_fd_sc_hd__dfrtp_1
X_10844_ net974 _05576_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__nand2_1
XANTENNA__06575__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12874__Q final_design.data_from_mem\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13563_ clknet_leaf_156_clk _00794_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[551\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10775_ net75 net1055 vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12514_ _06176_ net358 net330 net1850 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13494_ clknet_leaf_128_clk _00725_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[482\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07653__A2 _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12445_ net1821 net209 net336 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__mux2_1
XANTENNA__08803__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12376_ net1587 net212 net271 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14115_ clknet_leaf_53_clk _01312_ net1159 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_11327_ net745 _03878_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14046_ clknet_leaf_48_clk _00007_ net1147 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11258_ net427 net574 _05959_ net315 net1757 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10209_ final_design.uart.BAUD_counter\[3\] _05093_ vssd1 vssd1 vccd1 vccd1 _05094_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_52_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11189_ net425 net568 _05898_ net315 net2219 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12465__A2 net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07420_ final_design.cpu.reg_window\[1\] final_design.cpu.reg_window\[33\] net931
+ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08516__S1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07351_ final_design.cpu.reg_window\[259\] final_design.cpu.reg_window\[291\] net943
+ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__mux2_1
XANTENNA__09094__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ final_design.cpu.reg_window\[582\] final_design.cpu.reg_window\[614\] net913
+ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09021_ _02067_ _02447_ net630 vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11728__A1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold201 final_design.cpu.reg_window\[728\] vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08205__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold212 final_design.cpu.reg_window\[963\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold223 final_design.cpu.reg_window\[730\] vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold234 final_design.cpu.reg_window\[844\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold245 final_design.cpu.reg_window\[211\] vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold256 final_design.cpu.reg_window\[172\] vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 final_design.cpu.reg_window\[973\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 final_design.cpu.reg_window\[838\] vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09923_ _04109_ _04398_ _04838_ _04222_ _04833_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_113_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout703 _01753_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_4
Xhold289 final_design.cpu.reg_window\[607\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout714 net716 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout725 net727 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__buf_4
XANTENNA_fanout397_A _06261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout736 net737 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__buf_2
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout747 net748 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_1
X_09854_ net477 _04406_ _04691_ net491 vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__a211o_1
XANTENNA__09544__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout758 net759 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1104_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09036__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ final_design.CPU_instr_adr\[23\] _01722_ vssd1 vssd1 vccd1 vccd1 _03756_
+ sky130_fd_sc_hd__and2_1
X_09785_ net96 _04179_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__xnor2_1
X_06997_ final_design.cpu.reg_window\[79\] final_design.cpu.reg_window\[111\] net907
+ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout564_A _06238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _01365_ _02064_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09857__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10467__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10467__B2 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11664__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ _01998_ _02061_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout731_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout829_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1094_X net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11154__X _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07618_ _02563_ _02568_ net729 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08598_ net891 _03542_ _03548_ _03535_ _03536_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_83_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07080__A _02030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07549_ _02496_ _02497_ _02498_ _02499_ net779 net792 vssd1 vssd1 vccd1 vccd1 _02500_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12129__C _05858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10560_ _05283_ _05303_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__nor2_1
XANTENNA__08832__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_130_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09219_ _03132_ _03162_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__and2b_1
X_14202__1271 vssd1 vssd1 vccd1 vccd1 _14202__1271/HI net1271 sky130_fd_sc_hd__conb_1
X_10491_ _04040_ _05237_ _05238_ _04042_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12230_ net232 net2265 net374 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__mux2_1
XANTENNA__09388__A2 _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06424__A final_design.data_from_mem\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06438__1 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout986_X net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11195__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12161_ net176 net2304 net385 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_145_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11112_ _05831_ _05830_ final_design.uart.bits_received\[0\] vssd1 vssd1 vccd1 vccd1
+ _00205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09735__A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12092_ net579 _06082_ net511 net393 net1621 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__a32o_1
Xhold790 final_design.cpu.reg_window\[139\] vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11476__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ _05765_ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__nor2_1
XANTENNA__08899__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12869__Q final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12994_ net1336 _00225_ net1159 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09470__A _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11945_ _06146_ net292 net411 net2392 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12100__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11876_ net2510 net522 _06245_ net435 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13615_ clknet_leaf_93_clk _00846_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[603\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11407__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10827_ net45 _05558_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12080__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13546_ clknet_leaf_1_clk _00777_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[534\]
+ sky130_fd_sc_hd__dfrtp_1
X_10758_ net974 _05494_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13477_ clknet_leaf_17_clk _00708_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[465\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10689_ _05427_ _05428_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_97_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12428_ _06115_ net350 net340 net2312 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12383__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12359_ net2350 net362 net356 _06068_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__a22o_1
XANTENNA__07864__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07717__X _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06920_ final_design.cpu.reg_window\[978\] final_design.cpu.reg_window\[1010\] net903
+ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__mux2_1
X_14029_ clknet_leaf_139_clk _01260_ net1181 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1017\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11894__A0 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ net772 _01801_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__nor2_1
XANTENNA__09551__A2 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06996__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09570_ net559 net558 net556 net555 net455 net464 vssd1 vssd1 vccd1 vccd1 _04489_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_160_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06782_ final_design.cpu.reg_window\[22\] final_design.cpu.reg_window\[54\] net902
+ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__mux2_1
X_08521_ final_design.cpu.reg_window\[962\] final_design.cpu.reg_window\[994\] net865
+ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11646__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10449__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08708__B _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08452_ net722 _03396_ net731 vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09530__D _04448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07403_ _02350_ _02351_ _02352_ _02353_ net785 net794 vssd1 vssd1 vccd1 vccd1 _02354_
+ sky130_fd_sc_hd__mux4_1
X_08383_ final_design.cpu.reg_window\[70\] final_design.cpu.reg_window\[102\] net831
+ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07334_ final_design.cpu.reg_window\[964\] final_design.cpu.reg_window\[996\] net939
+ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__mux2_1
XANTENNA__12071__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07173__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10465__S net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07265_ final_design.cpu.reg_window\[326\] final_design.cpu.reg_window\[358\] net914
+ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout312_A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11788__C net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_A _01371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ _03683_ _03737_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07196_ _02143_ _02144_ _02145_ _02146_ net780 net799 vssd1 vssd1 vccd1 vccd1 _02147_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11177__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10385__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__A2 _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout500 _06264_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout779_A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 net512 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout522 net523 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_8
X_09906_ _04072_ _04824_ _04810_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_158_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout533 _02294_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_2
Xfanout544 _02026_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_2
Xfanout566 net568 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_2
X_09837_ net487 _04755_ _04341_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__a21o_1
XANTENNA__09542__A2 _04366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout577 net582 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__buf_2
Xfanout588 net597 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_2
XANTENNA__07553__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout599 net600 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout946_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ net321 _04683_ _04684_ net320 _04686_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08719_ _03669_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09699_ net547 net546 net545 net544 net454 net462 vssd1 vssd1 vccd1 vccd1 _04618_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11730_ net437 net592 _06223_ net298 net1917 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__a32o_1
XFILLER_0_166_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07014__S net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ net182 net641 vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ clknet_leaf_137_clk _00631_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[388\]
+ sky130_fd_sc_hd__dfrtp_1
X_10612_ _05354_ _05355_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_25_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11592_ net184 net645 vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13331_ clknet_leaf_31_clk _00562_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[319\]
+ sky130_fd_sc_hd__dfrtp_1
X_10543_ net94 final_design.VGA_adr\[2\] _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input75_A memory_size[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13262_ clknet_leaf_115_clk _00493_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[250\]
+ sky130_fd_sc_hd__dfrtp_1
X_10474_ net813 _05224_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12213_ net594 _06141_ net518 net379 net1581 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__a32o_1
X_13193_ clknet_leaf_95_clk _00424_ net1226 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[181\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10376__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12144_ net208 net2485 net385 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12075_ net575 _05959_ net509 net392 net1652 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__a32o_1
XANTENNA__10404__A _03450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ _05729_ _05733_ _05749_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06978__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2__f_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11628__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12977_ clknet_leaf_69_clk _00002_ net1244 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.current_client\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11928_ _06130_ net279 net408 net1892 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_72_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10851__A1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11859_ net2371 net521 _06241_ net430 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06616__X _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07155__S0 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13529_ clknet_leaf_166_clk _00760_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[517\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_166_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07050_ _01996_ _02000_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__clkbuf_4
XANTENNA__09221__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_81_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09375__A _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07952_ _02838_ _02901_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__nand2_1
XANTENNA__12659__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07619__A1_N net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06903_ _01853_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__inv_2
XANTENNA_wire535_X net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11867__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07883_ net552 _02832_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__nand2b_2
X_09622_ _02868_ net446 net443 _02866_ _04535_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__o221ai_1
XANTENNA__09822__B _04153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06834_ net900 _01777_ _01783_ _01765_ _01771_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a32o_2
X_14201__1270 vssd1 vssd1 vccd1 vccd1 _14201__1270/HI net1270 sky130_fd_sc_hd__conb_1
XANTENNA__11882__A3 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07623__A _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _02935_ _04471_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06765_ net767 _01715_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_108_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08504_ _02325_ net494 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_90_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12292__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__S1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09484_ _04401_ _04402_ net476 vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06696_ final_design.cpu.reg_window\[985\] final_design.cpu.reg_window\[1017\] net940
+ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__mux2_1
XANTENNA__09693__D1 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ net611 _03384_ _03360_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1171_A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07769__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ final_design.cpu.reg_window\[583\] final_design.cpu.reg_window\[615\] net833
+ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__mux2_1
XANTENNA__11799__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11398__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12972__Q final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12595__B2 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07317_ net535 _02267_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08297_ final_design.cpu.reg_window\[649\] final_design.cpu.reg_window\[681\] net842
+ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__mux2_1
XANTENNA__07697__S1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10070__A2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07248_ net759 _02198_ net754 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout896_A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10358__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ _02127_ _02128_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07449__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1224_X net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10190_ _05066_ _05079_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__nand2_4
XFILLER_0_44_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout330 _06284_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_4
Xfanout341 net342 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_8
Xfanout352 _06277_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09515__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout363 _06276_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_4
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_8
Xfanout385 _06266_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_6
X_12900_ clknet_leaf_68_clk _00138_ net1221 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11754__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_6
X_13880_ clknet_leaf_138_clk _01111_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[868\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12831_ net1368 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12762_ _06397_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__inv_2
XANTENNA__12283__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10833__A1 _04571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11713_ net600 _06016_ net637 vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12693_ final_design.VGA_data_control.v_count\[6\] _01403_ vssd1 vssd1 vccd1 vccd1
+ _06334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11644_ net426 net570 _06179_ net299 net1598 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_42_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_942 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12882__Q final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12586__B2 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_11575_ net566 net420 _06143_ net303 net1714 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__a32o_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_94_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput38 mem_adr_start[11] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
X_13314_ clknet_leaf_20_clk _00545_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[302\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput49 mem_adr_start[21] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_4
X_10526_ _05270_ _05271_ _05272_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_131_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13245_ clknet_leaf_12_clk _00476_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[233\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10457_ net1510 net1048 _05212_ net248 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_90_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08370__Y _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11010__A1 _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13176_ clknet_leaf_131_clk _00407_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[164\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08303__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ _03648_ _04991_ _04987_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08962__B1 final_design.CPU_instr_adr\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _06094_ net518 vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__nand2_4
XFILLER_0_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11849__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ net1870 net176 net397 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__mux2_1
XANTENNA__11313__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ _05733_ _05734_ net1457 net1046 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07612__S1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06550_ final_design.reqhand.instruction\[31\] final_design.data_from_mem\[31\] net983
+ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__mux2_1
XANTENNA__12274__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10824__A1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10824__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06481_ final_design.cpu.reg_window\[30\] final_design.cpu.reg_window\[62\] net928
+ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08220_ final_design.cpu.reg_window\[459\] final_design.cpu.reg_window\[491\] net857
+ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08274__A _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08151_ _03099_ _03100_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08245__A2 _03192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07102_ final_design.cpu.reg_window\[652\] final_design.cpu.reg_window\[684\] net928
+ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
XANTENNA__09657__X _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08082_ _02965_ _02996_ _03028_ _03032_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__o31ai_4
XANTENNA__08650__C1 _01597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11839__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07033_ final_design.cpu.reg_window\[782\] final_design.cpu.reg_window\[814\] net925
+ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08721__B _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07177__X _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08984_ final_design.CPU_instr_adr\[17\] net1026 _03916_ _03920_ vssd1 vssd1 vccd1
+ vccd1 _00228_ sky130_fd_sc_hd__a22o_1
X_07935_ _02882_ _02883_ _02884_ _02885_ net682 net704 vssd1 vssd1 vccd1 vccd1 _02886_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout477_A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07866_ net728 _02816_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__nor2_1
XANTENNA__09044__S net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09605_ _04446_ _04523_ _04228_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__o21ai_1
X_06817_ final_design.cpu.reg_window\[469\] final_design.cpu.reg_window\[501\] net963
+ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__mux2_1
X_07797_ final_design.cpu.reg_window\[153\] final_design.cpu.reg_window\[185\] net870
+ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout644_A _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout265_X net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09536_ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__inv_2
XANTENNA__12265__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06748_ final_design.cpu.reg_window\[23\] final_design.cpu.reg_window\[55\] net925
+ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__mux2_1
XANTENNA__08469__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09467_ net85 _04192_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__nand2_1
X_06679_ net749 _01497_ net672 _01629_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__a211o_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout909_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12280__A3 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11162__X _05875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08418_ final_design.cpu.reg_window\[133\] final_design.cpu.reg_window\[165\] net821
+ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__mux2_1
XANTENNA__12017__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09398_ net482 _04302_ _04316_ _04109_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__a211o_1
XANTENNA__08184__A _02000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12418__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10028__C1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08349_ final_design.cpu.reg_window\[455\] final_design.cpu.reg_window\[487\] net834
+ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__mux2_1
XANTENNA__09433__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10043__A2 _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11240__A1 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11360_ final_design.data_from_mem\[26\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06049_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ _04999_ _05040_ _05164_ vssd1 vssd1 vccd1 vccd1 final_design.pixel_data sky130_fd_sc_hd__and3_1
XANTENNA__11749__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11791__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11291_ _04473_ net661 _05843_ _05988_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_46_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13030_ clknet_leaf_170_clk _00261_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10242_ final_design.uart.BAUD_counter\[15\] _05113_ net810 vssd1 vssd1 vccd1 vccd1
+ _05115_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08123__S net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08095__S1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11543__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07747__B2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ _05017_ _05061_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_state\[1\]
+ sky130_fd_sc_hd__nor2_1
Xfanout1103 net1104 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__buf_2
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1114 net1115 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_4
Xfanout1125 net1127 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__clkbuf_4
Xfanout1136 net1137 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input38_A mem_adr_start[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1148 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__clkbuf_4
Xfanout1158 net1164 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_137_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11484__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1169 net1173 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout182 net183 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
XFILLER_0_156_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13932_ clknet_leaf_122_clk _01163_ net1217 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[920\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout193 _06031_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_2
XFILLER_0_88_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07263__A _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12877__Q final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13863_ clknet_leaf_13_clk _01094_ net1100 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[851\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12814_ net1374 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12256__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13794_ clknet_leaf_14_clk _01025_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[782\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _06359_ _06379_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12271__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06486__A1 final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12008__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12676_ _06325_ net1435 net994 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_146_Left_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ net213 net640 vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11231__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ net216 net643 vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__and2_1
Xwire561 _01535_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08273__A1_N net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10585__A3 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 final_design.cpu.reg_window\[970\] vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11782__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10509_ _05256_ _05257_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__nor2_1
Xhold619 final_design.cpu.reg_window\[668\] vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11489_ net184 net2444 net310 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13228_ clknet_leaf_123_clk _00459_ net1191 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[216\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ clknet_leaf_7_clk _00390_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[147\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_155_Left_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07720_ net621 _02668_ _02669_ net560 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a211oi_2
XANTENNA__12495__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ net891 _02583_ _02589_ _02595_ _02601_ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__o32a_4
XTAP_TAPCELL_ROW_105_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06602_ net762 _01552_ net756 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07582_ net726 _02532_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_157_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09321_ net464 _04237_ _04238_ _04239_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__a31o_1
XFILLER_0_165_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06533_ _01474_ _01481_ _01482_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__nor3_4
XTAP_TAPCELL_ROW_122_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09663__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12262__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09252_ _04167_ _04170_ _02609_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__a21o_1
XANTENNA__07620__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06464_ net1053 net1006 _01414_ vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08203_ final_design.cpu.reg_window\[718\] final_design.cpu.reg_window\[750\] net853
+ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09183_ net623 _03549_ _03523_ _01567_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08134_ final_design.cpu.reg_window\[589\] final_design.cpu.reg_window\[621\] net832
+ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__mux2_1
XANTENNA__10025__A2 _04398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06951__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11773__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ final_design.cpu.reg_window\[722\] final_design.cpu.reg_window\[754\] net818
+ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1134_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07016_ net936 _01852_ _01821_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a21bo_2
XANTENNA__07348__A _02294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout594_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ _01884_ _02457_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout761_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ _01755_ net618 vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__or2_1
XANTENNA__12486__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10502__A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08898_ _03799_ _03843_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__or2_1
X_07849_ net607 _02797_ _02773_ net553 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__o211a_1
XANTENNA__13463__RESET_B net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__inv_2
XANTENNA__12238__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09519_ net493 _04437_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10791_ _05525_ _05526_ net108 net1041 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12253__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06468__A1 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12530_ _02328_ _06193_ _06260_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__or3_1
XFILLER_0_136_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06427__A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07022__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14239__1304 vssd1 vssd1 vccd1 vccd1 _14239__1304/HI net1304 sky130_fd_sc_hd__conb_1
XFILLER_0_35_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12461_ net1836 net181 net338 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14200_ net1269 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
X_11412_ net2047 net241 net313 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__mux2_1
XANTENNA__07957__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12410__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06861__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12392_ net1575 net182 net272 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14131_ clknet_leaf_76_clk final_design.vga.h_next_count\[0\] net1254 vssd1 vssd1
+ vccd1 vccd1 final_design.VGA_data_control.h_count\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11479__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11343_ net748 _03859_ _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14062_ clknet_leaf_46_clk _00024_ net1149 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11274_ net426 net569 _05973_ net315 net1799 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_37_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13013_ clknet_leaf_41_clk _00244_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10225_ final_design.uart.BAUD_counter\[9\] _05103_ vssd1 vssd1 vccd1 vccd1 _05104_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_37_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10156_ net1061 _05050_ _05045_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold5 final_design.cpu.reg_window\[16\] vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12477__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12103__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09192__B net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ _04999_ _05002_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__or2_1
XANTENNA__10412__A _03321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13915_ clknet_leaf_155_clk _01146_ net1115 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[903\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload3_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13846_ clknet_leaf_125_clk _01077_ net1191 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[834\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13777_ clknet_leaf_108_clk _01008_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[765\]
+ sky130_fd_sc_hd__dfrtp_1
X_10989_ _01360_ _03844_ net1072 vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__mux2_1
XANTENNA__12244__A3 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11243__A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12728_ _06363_ _06361_ final_design.VGA_data_control.v_count\[1\] vssd1 vssd1 vccd1
+ vccd1 _06369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12659_ final_design.VGA_data_control.ready_data\[17\] net1032 net987 final_design.data_from_mem\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11204__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12401__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold405 final_design.cpu.reg_window\[50\] vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 final_design.cpu.reg_window\[764\] vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 final_design.cpu.reg_window\[754\] vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold438 final_design.cpu.reg_window\[58\] vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07168__A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold449 final_design.cpu.reg_window\[727\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09654__Y _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout907 net909 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_4
X_09870_ _03520_ _03521_ _03554_ _03555_ _04046_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__o311a_1
Xfanout918 net922 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_74_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 net933 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _03666_ _03771_ _03667_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a21o_1
XANTENNA__12180__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 final_design.cpu.reg_window\[291\] vssd1 vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07592__C1 _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1116 final_design.cpu.reg_window\[625\] vssd1 vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ final_design.CPU_instr_adr\[5\] net675 _01659_ vssd1 vssd1 vccd1 vccd1 _03703_
+ sky130_fd_sc_hd__and3_1
Xhold1127 final_design.cpu.reg_window\[303\] vssd1 vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12468__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1138 final_design.cpu.reg_window\[309\] vssd1 vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 final_design.reqhand.instruction\[20\] vssd1 vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07703_ _02650_ _02651_ _02652_ _02653_ net697 net715 vssd1 vssd1 vccd1 vccd1 _02654_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_124_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08683_ _03632_ _03633_ _02510_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07634_ final_design.cpu.reg_window\[28\] final_design.cpu.reg_window\[60\] net874
+ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06946__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ final_design.cpu.reg_window\[351\] final_design.cpu.reg_window\[383\] net844
+ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12235__A3 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09304_ net612 _03514_ _03516_ _02503_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_172_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06516_ net1051 net1008 net1005 final_design.reqhand.instruction\[3\] vssd1 vssd1
+ vccd1 vccd1 _01467_ sky130_fd_sc_hd__o31a_1
XFILLER_0_76_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ _02101_ _02446_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07111__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11994__A2 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09235_ _03326_ _03357_ _03324_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__a21oi_2
X_06447_ _01397_ _01400_ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__and2_1
XANTENNA__10992__A net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1251_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777__8 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__inv_2
XFILLER_0_118_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07777__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14009__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ _03419_ net488 vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08298__S1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08117_ net616 _03065_ _03066_ net543 vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11600__B net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09277__B net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09097_ _03711_ _03719_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1137_X net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08048_ final_design.cpu.reg_window\[466\] final_design.cpu.reg_window\[498\] net820
+ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__mux2_1
Xhold950 final_design.cpu.reg_window\[812\] vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold961 final_design.cpu.reg_window\[807\] vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold972 final_design.cpu.reg_window\[298\] vssd1 vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 final_design.cpu.reg_window\[931\] vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 final_design.cpu.reg_window\[641\] vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
X_10010_ _02326_ net455 _04238_ net468 vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__o211a_1
XANTENNA__06710__A _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ net452 _04907_ _04916_ net733 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a211o_2
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ _06163_ net289 net406 net1832 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09875__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08222__S1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11762__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10912_ net676 _05627_ _05638_ net976 _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__o221a_1
X_13700_ clknet_leaf_94_clk _00931_ net1227 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[688\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11682__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07812__Y _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ net245 net2112 net275 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13631_ clknet_leaf_133_clk _00862_ net1166 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[619\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10843_ final_design.CPU_instr_adr\[19\] net1013 _05572_ net1066 vssd1 vssd1 vccd1
+ vccd1 _05576_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_80_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09627__A1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12226__A3 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13562_ clknet_leaf_162_clk _00793_ net1105 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[550\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12631__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10774_ net75 net1055 vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12513_ _06175_ net345 net327 net1851 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__a22o_1
XANTENNA__07733__S0 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11985__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13493_ clknet_leaf_26_clk _00724_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[481\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_160_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_160_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_137_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12444_ net2522 net212 net336 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11198__A0 final_design.data_from_mem\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06591__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12890__Q final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12375_ net1981 net214 net272 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14114_ clknet_leaf_53_clk net1513 net1152 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11326_ net667 _03874_ net739 vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14045_ clknet_leaf_48_clk _00037_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11257_ net654 net209 vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_128_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10208_ _05093_ net811 _05092_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__and3b_1
XFILLER_0_158_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06620__A _01567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11188_ net654 net223 vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_52_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11238__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ final_design.vga.h_current_state\[0\] final_design.VGA_data_control.h_count\[8\]
+ final_design.VGA_data_control.h_count\[9\] final_design.vga.h_current_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__or4b_1
XANTENNA__09490__X _04409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09931__A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11672__S net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12465__A3 _06268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06619__X _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__Y _05947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13829_ clknet_leaf_150_clk _01060_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[817\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12217__A3 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07350_ final_design.cpu.reg_window\[323\] final_design.cpu.reg_window\[355\] net943
+ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11976__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07281_ _02228_ _02229_ _02230_ _02231_ net777 net797 vssd1 vssd1 vccd1 vccd1 _02232_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_151_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_151_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09020_ net2565 net1026 _03948_ _03952_ vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__a22o_1
XANTENNA__07597__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14102__RESET_B net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11189__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold202 final_design.cpu.reg_window\[732\] vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold213 final_design.cpu.reg_window\[250\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold224 final_design.cpu.reg_window\[530\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 final_design.cpu.reg_window\[1004\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold246 final_design.cpu.reg_window\[153\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold257 final_design.cpu.reg_window\[217\] vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 final_design.cpu.reg_window\[574\] vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold279 final_design.reqhand.instruction\[29\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _04341_ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_113_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout704 net707 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__buf_4
Xfanout715 net716 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_4
Xfanout726 net727 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout737 net738 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_8
X_09853_ _04741_ _04771_ net451 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07626__A _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08221__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout748 _01490_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout292_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 net766 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__buf_4
XANTENNA__11148__A _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14238__1303 vssd1 vssd1 vccd1 vccd1 _14238__1303/HI net1303 sky130_fd_sc_hd__conb_1
X_08804_ final_design.CPU_instr_adr\[23\] _01722_ vssd1 vssd1 vccd1 vccd1 _03755_
+ sky130_fd_sc_hd__or2_1
X_09784_ _04657_ _04678_ _04679_ _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__and4_1
X_06996_ _01943_ _01944_ _01945_ _01946_ net775 net796 vssd1 vssd1 vccd1 vccd1 _01947_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09306__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ final_design.CPU_instr_adr\[13\] _02030_ vssd1 vssd1 vccd1 vccd1 _03686_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09841__A _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout178_X net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1205_A final_design.cpu.reg_window\[411\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _01487_ _03615_ _03616_ _02094_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__o22a_4
XANTENNA__11664__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07617_ _02564_ _02565_ _02566_ _02567_ net696 net715 vssd1 vssd1 vccd1 vccd1 _02568_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08597_ net728 _03547_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__or2_2
XANTENNA__12208__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11416__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ final_design.cpu.reg_window\[543\] final_design.cpu.reg_window\[575\] net927
+ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__mux2_1
XANTENNA__09085__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07715__S0 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11967__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07479_ _02364_ _02429_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_142_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_142_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_162_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09218_ _03068_ _03099_ _03100_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10490_ net1068 _05237_ net1014 net1031 vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_17_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06705__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_101_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07079__Y _02030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09149_ _04056_ _04067_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09388__A3 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ net179 net2507 net385 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout979_X net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ _05830_ net1065 vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__and2b_1
XANTENNA__11757__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09735__B _04639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12091_ net592 _06075_ net518 net395 net1827 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_9_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold780 final_design.cpu.reg_window\[951\] vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold791 final_design.cpu.reg_window\[448\] vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09545__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11042_ _05760_ _05764_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11058__A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07970__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10897__A _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ net1335 _00224_ net1159 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11944_ _06145_ net290 net410 net1960 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__a22o_1
XANTENNA__12885__Q final_design.data_from_mem\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11875_ net189 net564 vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10826_ _05559_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__inv_2
X_13614_ clknet_leaf_117_clk _00845_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[602\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11407__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11958__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10757_ final_design.CPU_instr_adr\[15\] net1013 _05490_ net1066 vssd1 vssd1 vccd1
+ vccd1 _05494_ sky130_fd_sc_hd__a2bb2o_1
X_13545_ clknet_leaf_85_clk _00776_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[533\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_133_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_45_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09198__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06834__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13476_ clknet_leaf_106_clk _00707_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[464\]
+ sky130_fd_sc_hd__dfrtp_1
X_10688_ net70 final_design.VGA_adr\[9\] _05426_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__or3_1
XFILLER_0_153_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07210__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10408__Y _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12427_ _06114_ net358 net342 net1999 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10918__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08131__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09926__A _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ net2402 net363 net359 _06061_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__a22o_1
XANTENNA__10394__A1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11591__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11309_ net2459 net315 net420 _06004_ vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__a22o_1
X_12289_ net584 _06219_ net514 net370 net2095 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08339__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14028_ clknet_leaf_122_clk _01259_ net1197 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1016\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06850_ _01797_ _01798_ _01799_ _01800_ net787 net803 vssd1 vssd1 vccd1 vccd1 _01801_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_101_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06996__S1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06781_ final_design.cpu.reg_window\[86\] final_design.cpu.reg_window\[118\] net902
+ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_160_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08520_ final_design.cpu.reg_window\[770\] final_design.cpu.reg_window\[802\] net866
+ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__mux2_1
XANTENNA__11646__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10449__A2 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08451_ net728 _03401_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_69_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ final_design.cpu.reg_window\[514\] final_design.cpu.reg_window\[546\] net946
+ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08382_ _03329_ _03330_ _03331_ _03332_ net685 net700 vssd1 vssd1 vccd1 vccd1 _03333_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07078__A1 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07333_ final_design.cpu.reg_window\[772\] final_design.cpu.reg_window\[804\] net941
+ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11949__A2 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_124_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07173__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10737__A1_N net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07264_ _02213_ _02214_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__and2b_1
XFILLER_0_144_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09003_ _02002_ _02450_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__and2_1
XANTENNA__07120__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12246__B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12783__14 clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_115_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07195_ final_design.cpu.reg_window\[905\] final_design.cpu.reg_window\[937\] net924
+ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout305_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout501 _06264_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout512 net513 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__buf_4
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ _04819_ _04821_ _04823_ _04820_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__or4b_1
Xfanout523 _06239_ vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_8
Xfanout534 net535 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout674_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11334__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_X net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout556 net557 vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_4
Xfanout567 net568 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__dlymetal6s2s_1
X_09836_ _04606_ _04711_ net471 vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__mux2_1
Xfanout578 net582 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__buf_2
XANTENNA__07790__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout589 net591 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09571__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ net493 _04685_ _04117_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__o21a_1
X_06979_ net765 _01929_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout841_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08189__S0 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08718_ final_design.CPU_instr_adr\[20\] _01823_ vssd1 vssd1 vccd1 vccd1 _03669_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09698_ _03100_ net441 net442 _03099_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08649_ _02769_ _03597_ _03598_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11660_ net592 net424 _06187_ net302 net1546 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__a32o_1
XFILLER_0_166_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10611_ _05334_ _05337_ _05353_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_25_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11591_ net589 net423 _06151_ net305 net1572 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_115_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13330_ clknet_leaf_27_clk _00561_ net1139 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[318\]
+ sky130_fd_sc_hd__dfrtp_1
X_10542_ net95 final_design.VGA_adr\[3\] vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__xor2_1
XANTENNA__11270__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13261_ clknet_leaf_139_clk _00492_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[249\]
+ sky130_fd_sc_hd__dfrtp_1
X_10473_ final_design.CPU_instr_adr\[1\] net79 net1068 vssd1 vssd1 vccd1 vccd1 _05224_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12212_ net569 _06140_ net506 net376 net1889 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13192_ clknet_leaf_118_clk _00423_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[180\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input68_A memory_size[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10376__B2 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11487__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12143_ net209 net2253 net384 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12074_ net579 _05952_ net511 net393 net1463 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__a32o_1
XANTENNA__10404__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ _05729_ _05733_ _05749_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11876__B2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06978__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11628__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ clknet_leaf_73_clk _00001_ net1244 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.current_client\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11927_ net2513 net410 _06253_ net432 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ net212 net563 vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_99_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10809_ _05522_ _05540_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12053__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_106_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11789_ net2452 net413 _06233_ net430 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07155__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13528_ clknet_leaf_131_clk _00759_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[516\]
+ sky130_fd_sc_hd__dfrtp_1
X_14237__1302 vssd1 vssd1 vccd1 vccd1 _14237__1302/HI net1302 sky130_fd_sc_hd__conb_1
XFILLER_0_125_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11800__B2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13459_ clknet_leaf_31_clk _00690_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[447\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07875__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12356__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10367__B2 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_140_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07783__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ _02838_ _02901_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_162_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06902_ net754 net671 _01821_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__o21ai_4
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ net618 _02830_ _02831_ net552 vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__a211oi_1
X_06833_ net900 _01777_ _01783_ _01765_ _01771_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__a32oi_4
XANTENNA_wire528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ _04342_ _04539_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__and2b_1
X_09552_ _03590_ _04143_ _04157_ _03587_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__o31a_1
X_06764_ _01711_ _01712_ _01713_ _01714_ net776 net791 vssd1 vssd1 vccd1 vccd1 _01715_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_108_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08503_ net625 _03450_ _03451_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09483_ net547 net546 net545 net544 net457 net466 vssd1 vssd1 vccd1 vccd1 _04402_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06695_ final_design.cpu.reg_window\[793\] final_design.cpu.reg_window\[825\] net947
+ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09693__C1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_144_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08434_ _02267_ net611 vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__and2_1
XANTENNA__06954__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08365_ final_design.cpu.reg_window\[647\] final_design.cpu.reg_window\[679\] net856
+ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11799__C net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1164_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ net675 _01659_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08296_ final_design.cpu.reg_window\[713\] final_design.cpu.reg_window\[745\] net842
+ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_159_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07247_ _02194_ _02195_ _02196_ _02197_ net778 net797 vssd1 vssd1 vccd1 vccd1 _02198_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout210_X net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12347__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09748__B1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06542__X _01493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07178_ _02127_ _02128_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout791_A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08470__A _02294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10358__B2 final_design.data_from_mem\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout889_A net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1217_X net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout320 _04084_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout331 net332 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout342 _06279_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_8
Xfanout353 net354 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09515__A3 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout364 net365 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_6
Xfanout375 _06272_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_8
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_8
X_09819_ _03294_ _03569_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__nand2_1
Xfanout397 _06261_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_6
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12830_ net1370 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07025__S net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12761_ _06339_ _06391_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__or2_1
XANTENNA__08487__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11712_ net435 net587 _06214_ net297 net1616 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__a32o_1
X_12692_ _05008_ net967 _05059_ net808 net2563 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__a32o_1
XANTENNA__10833__A2 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12035__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11643_ net199 net638 vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10046__B1 _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08334__S0 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11574_ net201 net642 vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_1
XFILLER_0_135_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 mem_adr_start[12] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
X_10525_ _05270_ _05271_ _05272_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__and3_1
X_13313_ clknet_leaf_151_clk _00544_ net1116 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[301\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12338__A2 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ clknet_leaf_147_clk _00475_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[232\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10456_ _02602_ net602 vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11010__A2 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ clknet_leaf_145_clk _00406_ net1183 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[163\]
+ sky130_fd_sc_hd__dfrtp_1
X_10387_ net1378 net1045 _05174_ vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12106__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10415__A _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ net1642 net176 net389 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__mux2_1
XANTENNA__06973__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ net1841 net178 net397 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11008_ _05711_ _05731_ _05732_ net1018 vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__a31o_1
XANTENNA__12510__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07073__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11077__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12274__A1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ clknet_leaf_57_clk _00197_ net1162 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06480_ final_design.cpu.reg_window\[94\] final_design.cpu.reg_window\[126\] net929
+ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__mux2_1
XANTENNA__08555__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08150_ _03099_ _03100_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__nor2_1
XANTENNA__09978__B1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07101_ final_design.cpu.reg_window\[716\] final_design.cpu.reg_window\[748\] net928
+ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08081_ net550 _02996_ _03024_ _02993_ net551 vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__o32a_1
XFILLER_0_99_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13510__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07032_ final_design.cpu.reg_window\[846\] final_design.cpu.reg_window\[878\] net925
+ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__mux2_1
XANTENNA__06803__A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07205__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ net257 _03918_ net1026 vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07934_ final_design.cpu.reg_window\[918\] final_design.cpu.reg_window\[950\] net822
+ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__mux2_1
XANTENNA__09833__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06949__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12501__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07865_ _02812_ _02813_ _02814_ _02815_ net695 net712 vssd1 vssd1 vccd1 vccd1 _02816_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10512__A1 final_design.CPU_instr_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10512__B2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout372_A net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09604_ net487 _04437_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__nand2_1
XANTENNA__08181__A2 _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06816_ final_design.cpu.reg_window\[277\] final_design.cpu.reg_window\[309\] net964
+ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07796_ final_design.cpu.reg_window\[217\] final_design.cpu.reg_window\[249\] net870
+ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09535_ _04188_ _04453_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_27_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06747_ final_design.cpu.reg_window\[87\] final_design.cpu.reg_window\[119\] net925
+ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout258_X net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout637_A _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11443__X _06094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09466_ _04382_ _04383_ net738 _04381_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06678_ net753 _01628_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__and2_1
XANTENNA__06684__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08465__A _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12983__Q final_design.CPU_instr_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08417_ final_design.cpu.reg_window\[197\] final_design.cpu.reg_window\[229\] net821
+ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09397_ net465 _04080_ _04315_ net474 vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__o211a_1
XFILLER_0_171_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12783__14_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout804_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ final_design.cpu.reg_window\[263\] final_design.cpu.reg_window\[295\] net834
+ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__mux2_1
XANTENNA__09848__X _04767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09969__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11776__B1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08279_ _03229_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__inv_2
X_10310_ net1061 final_design.VGA_data_control.h_count\[5\] _05153_ _05163_ vssd1
+ vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__a31o_1
X_11290_ net651 _05984_ _05987_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10241_ final_design.uart.BAUD_counter\[15\] _05113_ vssd1 vssd1 vccd1 vccd1 _05114_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10553__A1_N net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09292__S1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__A3 _06127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _05061_ _05063_ final_design.h_out vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_state\[0\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10751__A1 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1104 net1164 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_4
Xfanout1115 net1118 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11765__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1126 net1127 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06859__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1137 net1156 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_2
Xfanout1148 net1149 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1159 net1160 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07544__A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13931_ clknet_leaf_15_clk _01162_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[919\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout183 _06067_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_2
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__buf_2
X_14236__1301 vssd1 vssd1 vccd1 vccd1 _14236__1301/HI net1301 sky130_fd_sc_hd__conb_1
XANTENNA__11700__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13862_ clknet_leaf_168_clk _01093_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[850\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12813_ net1451 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12256__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13793_ clknet_leaf_155_clk _01024_ net1113 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[781\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _05059_ _06373_ net967 vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__o21a_1
XANTENNA__06594__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12893__Q final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ final_design.VGA_data_control.ready_data\[25\] net1035 net990 final_design.data_from_mem\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input90_X net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12559__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09758__X _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ net431 net576 _06170_ net299 net1464 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__a32o_1
XANTENNA__08662__X _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11767__A0 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11231__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11557_ net577 net422 _06134_ net304 net1647 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__a32o_1
Xwire562 _01452_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10508_ final_design.CPU_instr_adr\[2\] net1073 final_design.CPU_instr_adr\[3\] vssd1
+ vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold609 final_design.cpu.reg_window\[278\] vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08314__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11488_ net185 net647 vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13227_ clknet_leaf_15_clk _00458_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[215\]
+ sky130_fd_sc_hd__dfrtp_1
X_10439_ net1389 net1040 _05203_ net246 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13158_ clknet_leaf_171_clk _00389_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[146\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12903__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12109_ net1866 net208 net389 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__mux2_1
X_13089_ clknet_leaf_159_clk _00320_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08148__C1 _02026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11298__A2 _05994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12495__A1 _06155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ net728 _02600_ net891 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_105_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06601_ _01548_ _01549_ _01550_ _01551_ net786 net804 vssd1 vssd1 vccd1 vccd1 _01552_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12247__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ _02528_ _02529_ _02530_ _02531_ net687 net708 vssd1 vssd1 vccd1 vccd1 _02532_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_157_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09320_ net464 _03639_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__nor2_1
X_06532_ _01478_ _01479_ _01457_ _01459_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_122_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13762__RESET_B net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09251_ _02673_ _02705_ _04168_ _04169_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__o31a_1
XFILLER_0_29_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06463_ _01405_ _01412_ _00211_ vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_174_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08202_ net719 _03152_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_174_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ _04097_ _04099_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__nor2_1
XANTENNA__13009__RESET_B net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11758__A0 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08133_ net718 _03077_ net730 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10754__S net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12094__X _06265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09820__C1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout218_A _05928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_6__f_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_71_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08064_ _03011_ _03012_ _03013_ _03014_ net682 net704 vssd1 vssd1 vccd1 vccd1 _03015_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08224__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10981__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ _01953_ _01954_ _01965_ net894 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_102_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07348__B _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_4__f_clk_X clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1127_A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout587_A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ final_design.CPU_instr_adr\[19\] net1049 _03904_ vssd1 vssd1 vccd1 vccd1
+ _00230_ sky130_fd_sc_hd__o21a_1
XANTENNA__11289__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07917_ _02866_ _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__or2_2
X_08897_ final_design.CPU_instr_adr\[26\] _03798_ vssd1 vssd1 vccd1 vccd1 _03843_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout754_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08179__B _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_95_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07848_ net607 _02797_ _02773_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07651__X _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12238__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ _02724_ _02729_ net721 vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ _04204_ _04336_ net475 vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__mux2_1
X_10790_ _05508_ _05524_ net1018 vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12429__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11997__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09449_ _04296_ _04364_ net474 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12460_ net1776 net182 net337 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__mux2_1
XANTENNA__08923__A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11749__A0 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11411_ net2012 net229 net312 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__mux2_1
X_12391_ net2031 net185 net273 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14130_ clknet_leaf_74_clk final_design.vga.v_next_state\[1\] net1246 vssd1 vssd1
+ vccd1 vccd1 final_design.vga.v_current_state\[1\] sky130_fd_sc_hd__dfrtp_1
X_11342_ net670 _03857_ net745 vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14061_ clknet_leaf_46_clk _00023_ net1149 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11273_ net654 net206 vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input50_A mem_adr_start[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _05103_ net811 _05102_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_37_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13012_ clknet_leaf_102_clk _00243_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11495__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10155_ _05045_ _05051_ _05052_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[3\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_89_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12888__Q final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10086_ _01369_ _01397_ _01398_ _05001_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__and4_1
Xhold6 final_design.cpu.reg_window\[26\] vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10412__B _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_86_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ clknet_leaf_163_clk _01145_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[902\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13845_ clknet_leaf_24_clk _01076_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[833\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08528__S0 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11524__A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15__f_clk_X clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13776_ clknet_leaf_115_clk _01007_ net1204 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[764\]
+ sky130_fd_sc_hd__dfrtp_1
X_10988_ _04529_ net252 vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__nor2_1
XANTENNA__06618__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11988__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12727_ final_design.VGA_data_control.v_count\[1\] _06361_ _06363_ _06367_ vssd1
+ vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12658_ _06316_ net1494 net991 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07408__A1 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10574__S net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11609_ net241 net640 vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12589_ net1530 net1011 net997 final_design.data_from_mem\[7\] vssd1 vssd1 vccd1
+ vccd1 _01282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_10_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08081__B2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold406 final_design.cpu.reg_window\[228\] vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 final_design.cpu.reg_window\[788\] vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold428 final_design.cpu.reg_window\[128\] vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold439 final_design.cpu.reg_window\[649\] vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10715__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__A0 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 net909 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10715__B2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout919 net922 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _03768_ _03769_ _03668_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_74_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_14__f_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
Xhold1106 final_design.cpu.reg_window\[51\] vssd1 vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 final_design.cpu.reg_window\[736\] vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _03700_ _03701_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__and2_1
Xhold1128 final_design.cpu.reg_window\[891\] vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_77_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1139 final_design.cpu.reg_window\[815\] vssd1 vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07702_ final_design.cpu.reg_window\[155\] final_design.cpu.reg_window\[187\] net881
+ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07344__A0 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08682_ _03611_ _03630_ _03628_ _03612_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07633_ final_design.cpu.reg_window\[92\] final_design.cpu.reg_window\[124\] net874
+ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07564_ _02504_ net612 vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__nand2_1
XANTENNA__08219__S net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11979__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06515_ final_design.data_from_mem\[3\] net1053 net1006 net1003 vssd1 vssd1 vccd1
+ vccd1 _01466_ sky130_fd_sc_hd__and4_1
X_09303_ net603 _04219_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_172_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07495_ _02130_ _02159_ _02443_ _02129_ _02099_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__o311a_1
XFILLER_0_119_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout335_A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1077_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06446_ final_design.VGA_data_control.v_count\[7\] final_design.VGA_data_control.v_count\[8\]
+ final_design.VGA_data_control.v_count\[5\] final_design.VGA_data_control.v_count\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__or4_2
XFILLER_0_17_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ _03390_ _03423_ _04148_ _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__a31o_2
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09165_ net498 net490 vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout502_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1244_A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14235__1300 vssd1 vssd1 vccd1 vccd1 _14235__1300/HI net1300 sky130_fd_sc_hd__conb_1
X_08116_ net616 _03065_ _03066_ net543 vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_16_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09096_ _02332_ _02431_ net632 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08047_ _01881_ net606 vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1032_X net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12156__A0 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold940 final_design.cpu.reg_window\[819\] vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold951 final_design.cpu.reg_window\[639\] vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 final_design.cpu.reg_window\[57\] vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09021__B1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07258__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold973 final_design.cpu.reg_window\[595\] vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 final_design.cpu.reg_window\[262\] vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold995 final_design.cpu.reg_window\[880\] vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout969_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10072__X _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11609__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10513__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ net452 _04907_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__a21o_1
X_08949_ _01825_ _02460_ net627 vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_32_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_68_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _06162_ net288 net406 net2156 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_174_Left_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10911_ _05639_ _05640_ net976 vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07430__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11682__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ net238 net2482 net275 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13630_ clknet_leaf_149_clk _00861_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[618\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10842_ net974 _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__or2_1
XANTENNA__09088__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789__20 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__inv_2
XFILLER_0_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13561_ clknet_leaf_166_clk _00792_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[549\]
+ sky130_fd_sc_hd__dfrtp_1
X_10773_ net251 _04697_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__and2b_1
XFILLER_0_55_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12631__B2 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07968__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07733__S1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12512_ _06174_ net351 net328 net1744 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__a22o_1
XANTENNA_input98_A memory_size[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13492_ clknet_leaf_141_clk _00723_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[480\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12443_ net2145 net214 net337 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11198__A1 final_design.reqhand.data_from_UART\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12374_ net1772 net215 net270 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__mux2_1
X_14113_ clknet_leaf_52_clk _01310_ net1159 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_105_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11325_ net438 net595 _06018_ net318 net1667 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14044_ clknet_leaf_49_clk _00036_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11256_ _04631_ net662 _05843_ _05957_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a211oi_4
XTAP_TAPCELL_ROW_128_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ final_design.uart.BAUD_counter\[1\] final_design.uart.BAUD_counter\[0\] final_design.uart.BAUD_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__and3_1
X_11187_ _04863_ net664 _05843_ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_52_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12114__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10423__A _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06620__B _01570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10138_ _01389_ final_design.vga.h_current_state\[1\] _05009_ vssd1 vssd1 vccd1 vccd1
+ _05040_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_59_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08118__A2 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10069_ _04987_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13828_ clknet_leaf_107_clk _01059_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[816\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13759_ clknet_leaf_135_clk _00990_ net1168 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[747\]
+ sky130_fd_sc_hd__dfrtp_1
X_07280_ final_design.cpu.reg_window\[902\] final_design.cpu.reg_window\[934\] net914
+ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06782__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11701__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11189__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10399__A1_N net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07179__A _02127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold203 final_design.cpu.reg_window\[978\] vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold214 final_design.VGA_data_control.ready_data\[0\] vssd1 vssd1 vccd1 vccd1 net1567
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold225 final_design.cpu.reg_window\[709\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__A0 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold236 final_design.cpu.reg_window\[778\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold247 final_design.cpu.reg_window\[212\] vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 net136 vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09921_ _04643_ _04839_ net484 vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__mux2_1
Xhold269 final_design.cpu.reg_window\[181\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout705 net707 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09554__A1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout716 _01752_ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout727 _01720_ vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_4
X_09852_ _04153_ _04154_ _03293_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__a21oi_1
Xfanout738 _01492_ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 _01477_ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_4
XANTENNA__11361__B2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08803_ final_design.CPU_instr_adr\[23\] _01722_ vssd1 vssd1 vccd1 vccd1 _03754_
+ sky130_fd_sc_hd__nor2_1
X_09783_ _04697_ _04699_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__xor2_1
XANTENNA__10052__B _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06995_ final_design.cpu.reg_window\[399\] final_design.cpu.reg_window\[431\] net907
+ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout285_A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ final_design.CPU_instr_adr\[13\] _02030_ vssd1 vssd1 vccd1 vccd1 _03685_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09857__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07868__A1 final_design.cpu.reg_window\[820\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _01999_ _02028_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__nor2_1
XANTENNA__11664__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout452_A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07616_ final_design.cpu.reg_window\[925\] final_design.cpu.reg_window\[957\] net883
+ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__mux2_1
X_08596_ _03543_ _03544_ _03545_ _03546_ net694 net702 vssd1 vssd1 vccd1 vccd1 _03547_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07547_ final_design.cpu.reg_window\[607\] final_design.cpu.reg_window\[639\] net927
+ vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12613__B2 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout717_A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10624__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07715__S1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07478_ _02426_ _02427_ _02395_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11611__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09217_ _03070_ _03101_ _03134_ _03164_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__and4_1
X_06429_ final_design.VGA_data_control.h_count\[3\] vssd1 vssd1 vccd1 vccd1 _01384_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11103__S net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09148_ _04059_ _04066_ net495 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09079_ final_design.CPU_instr_adr\[6\] net1029 _04004_ vssd1 vssd1 vccd1 vccd1 _00217_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11110_ net1065 _05078_ _05088_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07817__A net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12090_ net590 _06068_ net516 net394 net1954 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__a32o_1
XANTENNA__08412__S net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09735__C _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 final_design.cpu.reg_window\[285\] vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold781 final_design.cpu.reg_window\[399\] vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ _05764_ _05760_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__and2b_1
Xhold792 final_design.cpu.reg_window\[907\] vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11352__A1 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07028__S net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ net1334 _00223_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10897__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11104__B2 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08505__C1 _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07403__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ _06144_ net280 net408 net2209 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11874_ _06110_ net290 net522 net1926 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13613_ clknet_leaf_137_clk _00844_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[601\]
+ sky130_fd_sc_hd__dfrtp_1
X_10825_ net45 _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11407__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12604__B2 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13544_ clknet_leaf_126_clk _00775_ net1193 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[532\]
+ sky130_fd_sc_hd__dfrtp_1
X_10756_ net977 _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13475_ clknet_leaf_2_clk _00706_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[463\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12109__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10687_ net70 final_design.VGA_adr\[9\] _05426_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12426_ _06113_ net356 net341 net1986 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08131__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12357_ net2359 net362 net356 _06053_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06902__Y _01853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11591__A1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ net655 net569 net199 vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12288_ net586 _06218_ net515 net370 net2049 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__a32o_1
XANTENNA__06631__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08339__A2 _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11249__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14027_ clknet_leaf_18_clk _01258_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1015\]
+ sky130_fd_sc_hd__dfrtp_1
X_11239_ net2442 net317 _05942_ net432 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11343__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12540__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11536__X _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06780_ net758 _01730_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_160_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06770__A1 final_design.data_from_mem\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08450_ _03397_ _03398_ _03399_ _03400_ net691 net711 vssd1 vssd1 vccd1 vccd1 _03401_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08246__A_N net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07401_ final_design.cpu.reg_window\[578\] final_design.cpu.reg_window\[610\] net946
+ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
X_08381_ final_design.cpu.reg_window\[262\] final_design.cpu.reg_window\[294\] net831
+ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07332_ final_design.cpu.reg_window\[836\] final_design.cpu.reg_window\[868\] net941
+ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06806__A _01750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08293__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07401__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07263_ _02211_ _02212_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06525__B _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12359__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09002_ final_design.CPU_instr_adr\[15\] net1026 _03931_ _03936_ vssd1 vssd1 vccd1
+ vccd1 _00226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07194_ final_design.cpu.reg_window\[969\] final_design.cpu.reg_window\[1001\] net924
+ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout200_A _06003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08740__B _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08232__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout502 net504 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__buf_4
X_09904_ _04565_ _04822_ net496 vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__a21oi_1
Xfanout513 _06259_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout524 net527 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_6
XANTENNA__11334__A1 net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07538__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1207_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12531__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout546 _01966_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_2
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ net487 _04442_ _04515_ _04117_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a211o_1
Xfanout568 net572 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_4
Xfanout579 net580 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_2
XANTENNA_fanout288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06687__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ net480 _04055_ _04397_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__or3_1
X_06978_ _01925_ _01926_ _01927_ _01928_ net788 net806 vssd1 vssd1 vccd1 vccd1 _01929_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09063__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11098__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08717_ _01361_ _01690_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__nor2_1
XANTENNA__08189__S1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11606__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ net736 _04613_ _04615_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout834_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09160__C1 _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08502__A2 _03450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08648_ _02769_ _03597_ _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__o21a_1
XFILLER_0_166_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08579_ final_design.cpu.reg_window\[64\] final_design.cpu.reg_window\[96\] net862
+ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10610_ _05334_ _05337_ _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09299__A _02503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11590_ net186 net644 vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__and2_1
XFILLER_0_107_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10541_ net95 final_design.VGA_adr\[3\] vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13260_ clknet_leaf_123_clk _00491_ net1191 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[248\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout991_X net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10472_ net734 _04805_ net252 _04990_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12211_ net578 _06139_ net512 net377 net2016 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__a32o_1
XANTENNA__08569__A2 _03514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13191_ clknet_leaf_7_clk _00422_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[179\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10376__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11573__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12142_ net212 net2281 net385 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12073_ net2396 net394 net502 _05942_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__a22o_1
XANTENNA__11325__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12522__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ _05747_ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__and2_1
XANTENNA__11876__A2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07553__Y _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06597__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12896__Q final_design.data_from_mem\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12975_ clknet_leaf_69_clk _00000_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.current_client\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_99_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12999__RESET_B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11926_ net565 net240 net644 vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12928__RESET_B net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11857_ net2536 net522 _06240_ net432 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10808_ _05508_ _05542_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11788_ net655 net565 net208 vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07221__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10419__Y _05193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13527_ clknet_leaf_144_clk _00758_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[515\]
+ sky130_fd_sc_hd__dfrtp_1
X_10739_ net41 _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_136_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11800__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ clknet_leaf_27_clk _00689_ net1139 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[446\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09757__A1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12409_ _06241_ net501 net340 net2544 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__clkbuf_4
X_13389_ clknet_leaf_139_clk _00620_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[377\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07768__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13787__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08965__C1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09148__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07950_ _02866_ _02867_ _02897_ _02899_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_162_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12513__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07891__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06901_ _01468_ net744 net750 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a21o_1
X_07881_ net608 _02830_ _02805_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11867__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ _04100_ _04491_ net485 vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__mux2_1
X_06832_ net773 _01782_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__or2_1
XANTENNA__12302__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ _02964_ _04046_ _04351_ _04456_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__a41o_1
X_06763_ final_design.cpu.reg_window\[535\] final_design.cpu.reg_window\[567\] net911
+ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09142__C1 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08502_ net625 _03450_ _03451_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06694_ final_design.cpu.reg_window\[857\] final_design.cpu.reg_window\[889\] net947
+ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__mux2_1
X_09482_ net552 net551 net549 net548 net457 net466 vssd1 vssd1 vccd1 vccd1 _04401_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08433_ _03371_ _03372_ _03383_ net888 vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_93_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08735__B _02030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08364_ final_design.cpu.reg_window\[711\] final_design.cpu.reg_window\[743\] net833
+ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07131__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11252__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ _02248_ _02254_ _02265_ net894 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_116_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08295_ final_design.cpu.reg_window\[521\] final_design.cpu.reg_window\[553\] net841
+ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout415_A _06227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1157_A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07246_ final_design.cpu.reg_window\[391\] final_design.cpu.reg_window\[423\] net916
+ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07177_ net749 _01505_ net674 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_4
XFILLER_0_42_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10358__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08470__B net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07367__A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout784_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout310 _06095_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12504__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout321 _04073_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout332 net334 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_8
Xfanout343 net346 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_4
Xfanout354 net357 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_2
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout951_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout365 net367 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__buf_6
Xfanout376 net377 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11617__A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout387 _06266_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_4
X_09818_ _04222_ _04726_ _04731_ _04736_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__o211a_1
XANTENNA__10521__A _04847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout398 net399 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09749_ _03195_ net442 net439 _03197_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12760_ _06339_ _06391_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__nand2_1
XANTENNA__08487__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11711_ net198 net636 vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12691_ _01390_ net967 net808 net2569 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11642_ net425 net566 _06178_ net299 net1492 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10046__A1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07041__S net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08334__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11573_ net571 net420 _06142_ net303 net1905 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07998__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input80_A memory_size[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13312_ clknet_leaf_35_clk _00543_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[300\]
+ sky130_fd_sc_hd__dfrtp_1
X_10524_ _05235_ _05252_ _05251_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__o21ai_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire766 _01427_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__buf_4
XFILLER_0_80_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13243_ clknet_leaf_155_clk _00474_ net1112 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[231\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10455_ net1521 net1047 _05211_ net248 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_131_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09203__A3 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ clknet_leaf_130_clk _00405_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[162\]
+ sky130_fd_sc_hd__dfrtp_1
X_10386_ wb_manage.curr_state\[1\] net1 wb_manage.curr_state\[2\] vssd1 vssd1 vccd1
+ vccd1 _05174_ sky130_fd_sc_hd__or3b_1
XFILLER_0_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10415__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12125_ net1835 net178 net389 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__mux2_1
XANTENNA__06973__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ net2248 net180 net399 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__mux2_1
XANTENNA__11849__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _05711_ _05732_ _05731_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12122__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10431__A _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07073__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ clknet_leaf_50_clk _00196_ net1155 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11482__A0 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07686__C1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11909_ final_design.cpu.reg_window\[407\] _05845_ vssd1 vssd1 vccd1 vccd1 _06249_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_138_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ clknet_leaf_71_clk _00127_ net1240 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_103_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07100_ net761 _02050_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11785__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08080_ net550 _03024_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__nor2_1
XANTENNA__06790__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07031_ net760 _01975_ net755 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__o21a_1
XFILLER_0_141_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10606__A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06803__B net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08982_ _03918_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07933_ final_design.cpu.reg_window\[982\] final_design.cpu.reg_window\[1014\] net822
+ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__mux2_1
XANTENNA__08166__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout198_A _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12032__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ final_design.cpu.reg_window\[148\] final_design.cpu.reg_window\[180\] net866
+ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__mux2_1
XANTENNA__10512__A2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ _02702_ net440 _04519_ _04521_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_127_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06815_ final_design.cpu.reg_window\[341\] final_design.cpu.reg_window\[373\] net963
+ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07795_ final_design.cpu.reg_window\[25\] final_design.cpu.reg_window\[57\] net870
+ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout365_A net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ net76 _04187_ net77 vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_27_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06746_ _01693_ _01694_ _01695_ _01696_ net781 net801 vssd1 vssd1 vccd1 vccd1 _01697_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__06965__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09465_ _04382_ _04383_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06677_ final_design.reqhand.instruction\[26\] final_design.data_from_mem\[26\] net986
+ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout532_A _02356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11172__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08416_ final_design.cpu.reg_window\[5\] final_design.cpu.reg_window\[37\] net821
+ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__mux2_1
XANTENNA__09418__A0 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12017__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ net469 _04104_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10028__A1 _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08347_ final_design.cpu.reg_window\[327\] final_design.cpu.reg_window\[359\] net834
+ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1062_X net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07796__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11056__C_N net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06553__X _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ _03227_ _03228_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__nor2_2
XFILLER_0_116_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout999_A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07229_ final_design.cpu.reg_window\[968\] final_design.cpu.reg_window\[1000\] net921
+ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10240_ _05113_ net810 _05112_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__and3b_1
XFILLER_0_132_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07827__S0 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ final_design.vga.h_current_state\[0\] final_design.vga.h_current_state\[1\]
+ _05016_ _05062_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__a31o_1
XANTENNA__09583__Y _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1105 net1111 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09516__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1116 net1117 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__clkbuf_4
Xfanout1127 net1128 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout954_X net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1138 net1145 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__clkbuf_4
Xfanout1149 net1156 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__clkbuf_2
X_13930_ clknet_leaf_165_clk _01161_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[918\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_35_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06707__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout184 _06060_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_2
Xfanout195 _06024_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_2
XANTENNA__11700__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13861_ clknet_leaf_150_clk _01092_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[849\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12812_ net1361 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__clkbuf_1
X_13792_ clknet_leaf_39_clk _01023_ net1136 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[780\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12743_ _05059_ _06373_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12674_ _06324_ net1442 net993 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__mux2_1
XANTENNA__12008__A2 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ net215 net638 vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_133_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07559__X _02510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input83_X net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11556_ net217 net643 vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__and2_1
XANTENNA__08632__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__A _01850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10507_ final_design.CPU_instr_adr\[3\] net1031 net1073 vssd1 vssd1 vccd1 vccd1 _05256_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_150_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12117__S net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11487_ net186 net2472 net309 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__mux2_1
XANTENNA__13308__RESET_B net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11519__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ clknet_leaf_0_clk _00457_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[214\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ _02991_ net601 vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12192__A1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13157_ clknet_leaf_5_clk _00388_ net1096 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[145\]
+ sky130_fd_sc_hd__dfrtp_1
X_10369_ net11 net1038 net1021 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1
+ vccd1 _00122_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_143_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ net1887 net209 net388 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__mux2_1
XANTENNA__08330__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13088_ clknet_leaf_36_clk _00319_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11257__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ net1635 net211 net397 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__mux2_1
XANTENNA__09896__A0 _02126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12495__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12943__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_158_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06600_ final_design.cpu.reg_window\[412\] final_design.cpu.reg_window\[444\] net955
+ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07580_ final_design.cpu.reg_window\[671\] final_design.cpu.reg_window\[703\] net846
+ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08566__A _02394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06531_ _01454_ _01455_ _01458_ _01460_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_122_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09250_ _02670_ _02702_ _02671_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__o21ba_1
X_06462_ _01405_ _01412_ _00211_ vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08201_ _03148_ _03149_ _03150_ _03151_ net688 net709 vssd1 vssd1 vccd1 vccd1 _03152_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_174_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08572__Y _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08132_ net727 _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_78_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06814__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ final_design.cpu.reg_window\[914\] final_design.cpu.reg_window\[946\] net818
+ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__mux2_1
XANTENNA__10430__B2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12027__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07014_ _01959_ _01964_ net759 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1022_A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ _03899_ _03900_ _03903_ net256 net1027 vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__a221o_1
XANTENNA__08240__S net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07916_ net618 _02863_ _02865_ net555 vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a211oi_2
XANTENNA__10071__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08234__S0 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08896_ _02471_ net632 _03839_ _03841_ net259 vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__a311o_1
XANTENNA__12486__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07847_ _01788_ net618 vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__nor2_1
XANTENNA__11694__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout270_X net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06695__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07778_ _02725_ _02726_ _02727_ _02728_ net695 net702 vssd1 vssd1 vccd1 vccd1 _02729_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09639__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07380__A _02326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09517_ net487 _04435_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06729_ final_design.cpu.reg_window\[600\] final_design.cpu.reg_window\[632\] net946
+ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout914_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09448_ net486 _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13819__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ net481 _04097_ _04296_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07379__X _02330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ net1712 net232 net314 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12390_ net1615 net187 net272 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__mux2_1
XANTENNA__12410__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11341_ net429 net578 _06032_ net316 net1783 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14060_ clknet_leaf_46_clk _00022_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11272_ _04509_ net662 _05843_ _05971_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_132_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13011_ net1353 _00242_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10223_ final_design.uart.BAUD_counter\[7\] final_design.uart.BAUD_counter\[8\] _05099_
+ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__and3_1
XANTENNA__08917__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input43_A mem_adr_start[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ _01384_ _05048_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_89_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10085_ final_design.VGA_data_control.v_count\[0\] _05000_ final_design.VGA_data_control.v_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12477__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 final_design.cpu.reg_window\[21\] vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_85_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913_ clknet_leaf_166_clk _01144_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[901\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13844_ clknet_leaf_105_clk _01075_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[832\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08528__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13775_ clknet_leaf_92_clk _01006_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[763\]
+ sky130_fd_sc_hd__dfrtp_1
X_10987_ _05710_ _05711_ _05713_ net1042 net1381 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__a32o_1
XANTENNA__06618__B _01568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12726_ final_design.VGA_data_control.v_count\[1\] _06366_ vssd1 vssd1 vccd1 vccd1
+ _06367_ sky130_fd_sc_hd__and2b_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07656__A2 _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12657_ final_design.VGA_data_control.ready_data\[16\] net1032 net987 final_design.data_from_mem\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08833__B final_design.CPU_instr_adr\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11608_ net2319 net300 _06161_ net428 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12588_ net2529 net1012 net998 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1
+ vccd1 _01281_ sky130_fd_sc_hd__a22o_1
XANTENNA__12401__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08325__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10427__Y _05197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11539_ net232 net2515 net305 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__mux2_1
Xhold407 final_design.cpu.reg_window\[702\] vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold418 final_design.cpu.reg_window\[441\] vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09945__A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold429 final_design.cpu.reg_window\[255\] vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12165__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13209_ clknet_leaf_168_clk _00440_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[197\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14189_ net1259 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_1_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout909 net912 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ final_design.CPU_instr_adr\[6\] _02240_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__or2_1
Xhold1107 net147 vssd1 vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1118 final_design.cpu.reg_window\[111\] vssd1 vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12468__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1129 final_design.cpu.reg_window\[390\] vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
X_07701_ final_design.cpu.reg_window\[219\] final_design.cpu.reg_window\[251\] net881
+ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08681_ _02545_ _03610_ _03631_ _02542_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_124_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08567__Y _03518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07471__Y _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ net721 _02582_ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__nor2_1
XANTENNA__12310__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07404__S net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07563_ _01488_ net746 net738 net670 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__or4_1
XFILLER_0_159_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09302_ net498 net603 _04111_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06514_ _01458_ _01460_ _01461_ _01462_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07494_ _02129_ _02444_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ _03324_ _04151_ _04150_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__o21ai_1
X_06445_ _01369_ _01398_ vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout230_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06950__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11450__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_A net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09164_ _04080_ _04082_ net469 vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__mux2_1
XANTENNA__08235__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06870__A3 _01495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08115_ _02064_ net616 vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__nor2_1
XANTENNA__10403__B2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10066__A _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09095_ net2549 net1030 _04018_ vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1237_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09855__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__or2_1
Xhold930 final_design.cpu.reg_window\[447\] vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold941 final_design.cpu.reg_window\[341\] vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold952 final_design.cpu.reg_window\[423\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap671 _01851_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_4
Xhold963 final_design.cpu.reg_window\[428\] vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07258__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold974 final_design.cpu.reg_window\[499\] vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 final_design.cpu.reg_window\[410\] vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 final_design.cpu.reg_window\[637\] vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11609__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14089__RESET_B net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ _04124_ _04915_ _04914_ _04911_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout864_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ final_design.CPU_instr_adr\[21\] _03888_ net1049 vssd1 vssd1 vccd1 vccd1
+ _00232_ sky130_fd_sc_hd__mux2_1
XANTENNA__08207__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09590__A _04502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08879_ net628 _03826_ _03824_ net260 vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a211o_1
XFILLER_0_169_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10910_ net1054 _05636_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__nor2_1
X_11890_ net224 net1934 net274 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__mux2_1
XANTENNA__07430__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07314__S net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10841_ net973 _05572_ _05573_ net968 vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_80_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09589__X _04508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12092__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13560_ clknet_leaf_129_clk _00791_ net1176 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[548\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ _05347_ _05385_ _05502_ _05507_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_149_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12631__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13653__RESET_B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12511_ _06173_ net347 net328 net1620 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13491_ clknet_leaf_32_clk _00722_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[479\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12442_ net1818 net215 net335 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12395__A1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12373_ net2140 net218 net271 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14112_ clknet_leaf_52_clk net1402 net1151 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11324_ net600 net658 net196 vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_56_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14043_ clknet_leaf_49_clk _00035_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11255_ net651 _05953_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11355__C1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10206_ final_design.uart.BAUD_counter\[1\] final_design.uart.BAUD_counter\[0\] final_design.uart.BAUD_counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_128_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11186_ net660 _05893_ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_52_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10423__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ net2560 net967 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.next_state\[1\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11658__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09946__S0 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10068_ _01495_ net253 _04044_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_141_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13827_ clknet_leaf_5_clk _01058_ net1096 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[815\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13758_ clknet_leaf_19_clk _00989_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[746\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12083__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08844__A final_design.CPU_instr_adr\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12709_ net1064 _06338_ _06343_ _06344_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__a22o_1
XANTENNA__06837__B1 _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11830__A0 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13689_ clknet_leaf_167_clk _00920_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[677\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11189__A2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12386__A1 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07179__B _02128_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold204 net121 vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold215 final_design.cpu.reg_window\[671\] vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold226 final_design.cpu.reg_window\[983\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold237 final_design.cpu.reg_window\[782\] vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09920_ _04778_ _04834_ net471 vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__mux2_1
Xhold248 final_design.cpu.reg_window\[490\] vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold259 final_design.cpu.reg_window\[700\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12305__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout706 net707 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_4
XFILLER_0_111_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09851_ _04181_ _04769_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout717 net718 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_4
XANTENNA__08211__C1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11897__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14182__RESET_B net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout728 net729 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 net742 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_2
X_08802_ _03670_ _03752_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__or2_1
XANTENNA__11361__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14111__RESET_B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09782_ _04697_ _04699_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06994_ final_design.cpu.reg_window\[463\] final_design.cpu.reg_window\[495\] net909
+ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__mux2_1
X_08733_ _03683_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout180_A _06074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09841__C _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12310__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08738__B _02097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout278_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ _02028_ _02061_ _03613_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__o21a_1
XANTENNA__12040__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07134__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07615_ final_design.cpu.reg_window\[989\] final_design.cpu.reg_window\[1021\] net880
+ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08595_ final_design.cpu.reg_window\[512\] final_design.cpu.reg_window\[544\] net871
+ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1187_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12074__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07546_ final_design.cpu.reg_window\[671\] final_design.cpu.reg_window\[703\] net927
+ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07477_ _02426_ _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout612_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11180__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _03589_ _04134_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__nand2_1
X_06428_ final_design.VGA_data_control.state\[0\] vssd1 vssd1 vccd1 vccd1 _01383_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_146_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12377__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09147_ _04060_ _04065_ net478 vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09078_ _03655_ _04002_ _04003_ net1050 vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11179__X _05890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08029_ final_design.cpu.reg_window\[787\] final_design.cpu.reg_window\[819\] net828
+ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__mux2_1
Xhold760 final_design.cpu.reg_window\[168\] vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11337__C1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold771 final_design.cpu.reg_window\[446\] vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold782 final_design.cpu.reg_window\[945\] vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ net88 _05737_ _05763_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__a21o_1
XANTENNA__11888__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09545__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold793 final_design.cpu.reg_window\[643\] vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__B1 final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07833__A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ net1333 _00222_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_11942_ _06143_ net278 net408 net2080 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07403__S1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11873_ net2252 net521 _06244_ net430 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13612_ clknet_leaf_125_clk _00843_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[600\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10824_ net676 _05546_ _05557_ net977 _05556_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__o221a_1
XANTENNA_input100_X net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12065__B1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06883__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06736__X _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07167__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13543_ clknet_leaf_10_clk _00774_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[531\]
+ sky130_fd_sc_hd__dfrtp_1
X_10755_ net973 _05490_ _05491_ _04042_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12080__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11090__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13474_ clknet_leaf_29_clk _00705_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[462\]
+ sky130_fd_sc_hd__dfrtp_1
X_10686_ net71 net1057 vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12425_ _06112_ net358 net342 net2481 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10379__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11040__A1 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12356_ net2545 net362 net355 _06046_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11307_ _04570_ net659 net598 _06002_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__o211a_2
XFILLER_0_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11591__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12125__S net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08419__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12287_ net572 _06217_ net507 net368 net1848 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__a32o_1
XANTENNA__10434__A _02929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14026_ clknet_leaf_3_clk _01257_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1014\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11249__B net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ net656 net583 net213 vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11879__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11169_ _05855_ _05880_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_143_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11265__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07400_ final_design.cpu.reg_window\[642\] final_design.cpu.reg_window\[674\] net946
+ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07889__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08380_ final_design.cpu.reg_window\[326\] final_design.cpu.reg_window\[358\] net831
+ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__mux2_1
XANTENNA__06646__X _01597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07331_ net764 _02275_ net756 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11803__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12071__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07262_ _02211_ _02212_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09001_ net630 _03934_ _03935_ net256 _03933_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__a311o_1
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07193_ final_design.cpu.reg_window\[777\] final_design.cpu.reg_window\[809\] net925
+ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07235__A0 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08513__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08983__B1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12035__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10790__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07129__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09903_ net488 _04559_ _04560_ _04262_ _04120_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__a221o_1
XANTENNA__11159__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout503 net504 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_2
XFILLER_0_10_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout514 net517 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout525 net527 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07538__A1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_A _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout536 _02239_ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12531__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout547 _01937_ vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_2
X_09834_ _03229_ _04087_ net441 _03227_ _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a221o_1
Xfanout569 net572 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__buf_2
X_09765_ _04393_ _04402_ net471 vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__mux2_1
XANTENNA__10888__A2_N _05615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06977_ final_design.cpu.reg_window\[912\] final_design.cpu.reg_window\[944\] net957
+ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout183_X net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11098__A1 _04177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ final_design.CPU_instr_adr\[25\] _01660_ vssd1 vssd1 vccd1 vccd1 _03667_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12295__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09696_ _01382_ _04185_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09160__B1 _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08647_ _01658_ _02765_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout827_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _03525_ _03526_ _03527_ _03528_ net692 net711 vssd1 vssd1 vccd1 vccd1 _03529_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12598__B2 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09999__C1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07529_ final_design.cpu.reg_window\[479\] final_design.cpu.reg_window\[511\] net933
+ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XANTENNA__09299__B net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10540_ net252 _04864_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__and2b_1
XANTENNA__11270__A1 _01967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10471_ net101 net1045 net1016 _05222_ vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12210_ net574 _06138_ net509 net376 net1562 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__a32o_1
X_13190_ clknet_leaf_171_clk _00421_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[178\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11573__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12141_ net213 net2410 net386 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07039__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12072_ net576 _05935_ net510 net392 net2098 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__a32o_1
Xhold590 final_design.cpu.reg_window\[89\] vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11325__A2 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ _05735_ _05746_ net55 vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__or3b_1
XFILLER_0_159_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06878__S net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11089__B2 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12974_ clknet_leaf_69_clk _00211_ net1244 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.current_client\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12286__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11925_ _06128_ net289 net410 net2036 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11372__X _06060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ net214 net564 vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ _05524_ _05540_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12589__B2 final_design.data_from_mem\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11787_ net2401 net412 net281 _05959_ vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10429__A _03129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10738_ net676 _05462_ _05475_ net977 _05474_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__o221a_1
X_13526_ clknet_leaf_130_clk _00757_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[514\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_41_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13457_ clknet_leaf_108_clk _00688_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[445\]
+ sky130_fd_sc_hd__dfrtp_1
X_10669_ _05408_ _05409_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12408_ _06240_ net502 net341 net2494 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__a22o_1
XANTENNA__12210__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ clknet_leaf_121_clk _00619_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[376\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08333__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12363__B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07768__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__clkbuf_4
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__clkbuf_4
X_12339_ _06231_ net502 net360 net2409 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__a22o_1
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06900_ _01468_ net743 net750 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a21oi_4
X_14009_ clknet_leaf_165_clk _01240_ net1083 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[997\]
+ sky130_fd_sc_hd__dfrtp_1
X_07880_ _01504_ _01822_ net608 vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__and3_1
XANTENNA__06788__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06831_ _01778_ _01779_ _01780_ _01781_ net789 net794 vssd1 vssd1 vccd1 vccd1 _01782_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11707__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ _04072_ _04468_ _04462_ _04464_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__or4b_1
XANTENNA__12277__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06762_ final_design.cpu.reg_window\[599\] final_design.cpu.reg_window\[631\] net911
+ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__mux2_1
XANTENNA__09142__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08501_ _02330_ net614 vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_108_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09481_ _04056_ _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06693_ net763 _01637_ net756 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12292__A3 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08432_ _03377_ _03382_ net717 vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08508__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08363_ _03310_ _03311_ _03312_ _03313_ net686 net706 vssd1 vssd1 vccd1 vccd1 _03314_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07314_ _02259_ _02264_ net758 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11252__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07456__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ final_design.cpu.reg_window\[585\] final_design.cpu.reg_window\[617\] net841
+ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07245_ final_design.cpu.reg_window\[455\] final_design.cpu.reg_window\[487\] net916
+ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout408_A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12201__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07176_ net895 _02119_ _02125_ _02107_ _02113_ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a32o_2
XFILLER_0_108_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12752__A1 final_design.VGA_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10074__A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout300 net302 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout311 net314 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_6
XANTENNA__11307__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 _04047_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_4
Xfanout333 net334 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_8
Xfanout344 net346 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_2
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09381__A0 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout366 net367 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_8
XANTENNA__11176__Y _05887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout377 _06271_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11617__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ _04378_ _04735_ net498 vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__a21o_1
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_6
XANTENNA__10521__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 _06261_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_4
XANTENNA__13426__RESET_B net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12268__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _04261_ _04262_ net496 _04097_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09679_ _04595_ _04596_ net737 _04594_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__o211ai_4
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12283__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ net570 net420 _06213_ net295 net1893 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__a32o_1
X_12690_ _01383_ final_design.VGA_data_control.state\[1\] _06332_ vssd1 vssd1 vccd1
+ vccd1 _06333_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07322__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11641_ net201 net638 vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09436__A1 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10046__A2 _04576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ net203 net642 vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_42_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13311_ clknet_leaf_137_clk _00542_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[299\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07998__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10523_ net94 final_design.VGA_adr\[2\] vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__or2_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11066__A1_N net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13242_ clknet_leaf_163_clk _00473_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[230\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input73_A memory_size[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ _02668_ net602 vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13173_ clknet_leaf_40_clk _00404_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[161\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10385_ net1596 net1041 net1015 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12124_ net1732 net180 net391 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12055_ net1628 net183 net398 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__mux2_1
X_11006_ net53 _05708_ _05712_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11019__S net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12259__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08676__X _03627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12957_ clknet_leaf_50_clk _00195_ net1155 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12274__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_116_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11908_ net816 _06246_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_138_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08328__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ clknet_leaf_87_clk _00126_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09013__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11839_ net182 net1910 net268 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08635__C1 _01938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11785__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13509_ clknet_leaf_17_clk _00740_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[497\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08650__A2 _02668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07030_ net769 _01980_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10606__B final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08938__B1 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12734__B2 final_design.VGA_data_control.v_count\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_141_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14219__1288 vssd1 vssd1 vccd1 vccd1 _14219__1288/HI net1288 sky130_fd_sc_hd__conb_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08981_ _03793_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__or2_2
XANTENNA__11277__X _05976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07932_ final_design.cpu.reg_window\[790\] final_design.cpu.reg_window\[822\] net822
+ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__mux2_1
XANTENNA__12498__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12313__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08166__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08299__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10843__A1_N final_design.CPU_instr_adr\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ final_design.cpu.reg_window\[212\] final_design.cpu.reg_window\[244\] net868
+ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__mux2_1
X_09602_ _04074_ _04440_ _04517_ net499 _04520_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__o221a_1
X_06814_ net773 _01764_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_127_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07794_ final_design.cpu.reg_window\[89\] final_design.cpu.reg_window\[121\] net870
+ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09533_ net737 _04429_ _04450_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__nand3_4
XFILLER_0_155_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06745_ final_design.cpu.reg_window\[407\] final_design.cpu.reg_window\[439\] net934
+ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout260_A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09666__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08469__A2 _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12265__A3 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ _02735_ _02769_ _04281_ net450 vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08238__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06676_ net898 _01619_ _01625_ _01612_ _01613_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__a32o_4
XFILLER_0_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08415_ final_design.cpu.reg_window\[69\] final_design.cpu.reg_window\[101\] net821
+ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__mux2_1
XANTENNA__11172__B net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09418__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09395_ _02576_ _04087_ net445 _02575_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_58_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout525_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11225__A1 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ _02212_ net618 vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__or2_1
XANTENNA__12422__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09969__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08762__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06834__X _01785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11776__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08277_ net604 _03224_ _03200_ net540 vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07228_ final_design.cpu.reg_window\[776\] final_design.cpu.reg_window\[808\] net942
+ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout894_A _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07159_ final_design.cpu.reg_window\[202\] final_design.cpu.reg_window\[234\] net934
+ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
XANTENNA__09051__C1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07827__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10170_ final_design.vga.h_current_state\[0\] _05009_ vssd1 vssd1 vccd1 vccd1 _05062_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1106 net1111 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_4
Xfanout1117 net1118 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12489__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1128 net1164 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__clkbuf_4
Xfanout1139 net1145 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_156_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout185 _06060_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13260__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout947_X net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 _06016_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11700__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13860_ clknet_leaf_106_clk _01091_ net1205 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[848\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09106__A0 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12811_ net1356 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__clkbuf_1
X_13791_ clknet_leaf_138_clk _01022_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[779\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12256__A3 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12742_ _06359_ _06379_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__or2_1
XANTENNA__07052__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12673_ final_design.VGA_data_control.ready_data\[24\] net1034 net989 final_design.data_from_mem\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07987__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ net577 net422 _06169_ net300 net1461 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__a32o_1
XANTENNA__11216__B2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12413__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11810__B net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11555_ net427 net575 _06133_ net303 net2113 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__a32o_1
Xwire531 _02389_ vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ _05235_ _05254_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_150_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11486_ net187 net647 vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_150_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13225_ clknet_leaf_85_clk _00456_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[213\]
+ sky130_fd_sc_hd__dfrtp_1
X_10437_ net255 _05202_ net1040 net1602 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_27_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13156_ clknet_leaf_94_clk _00387_ net1227 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[144\]
+ sky130_fd_sc_hd__dfrtp_1
X_10368_ net10 net1038 net1021 final_design.data_from_mem\[17\] vssd1 vssd1 vccd1
+ vccd1 _00121_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13348__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12107_ net1593 net211 net389 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__mux2_1
XANTENNA__11538__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ clknet_leaf_133_clk _00318_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12133__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10442__A _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10299_ _05149_ _05151_ _05152_ _01384_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__o22a_1
XANTENNA__07227__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12038_ net2198 net213 net398 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__mux2_1
XANTENNA__09896__A1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__B _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07751__A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13989_ clknet_leaf_150_clk _01220_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[977\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12247__A3 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11273__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06530_ _01478_ _01479_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__and2_2
XANTENNA__07470__B net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12983__RESET_B net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06461_ net1073 final_design.reqhand.current_client\[1\] _01393_ vssd1 vssd1 vccd1
+ vccd1 _00211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08200_ final_design.cpu.reg_window\[910\] final_design.cpu.reg_window\[942\] net843
+ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12404__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09180_ net481 _04098_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_174_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08131_ _03078_ _03079_ _03080_ _03081_ net685 net706 vssd1 vssd1 vccd1 vccd1 _03082_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12308__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09965__X _04884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08062_ final_design.cpu.reg_window\[978\] final_design.cpu.reg_window\[1010\] net820
+ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10430__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07013_ _01960_ _01961_ _01962_ _01963_ net775 net791 vssd1 vssd1 vccd1 vccd1 _01964_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08521__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11448__A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06493__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12043__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1015_A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ net607 _02863_ _02839_ net555 vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__o211a_1
X_08895_ net632 _03840_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__nor2_1
XANTENNA__09887__A1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08234__S1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11694__A1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ net893 _02796_ _02785_ _02784_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__09205__X _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ final_design.cpu.reg_window\[536\] final_design.cpu.reg_window\[568\] net865
+ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12238__A3 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_A _06123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07380__B _02330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06728_ _01675_ _01676_ _01677_ _01678_ net787 net793 vssd1 vssd1 vccd1 vccd1 _01679_
+ sky130_fd_sc_hd__mux4_1
X_09516_ _04337_ _04434_ net475 vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07745__S0 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11997__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09447_ net481 _04362_ _04363_ _04365_ _04293_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__o32a_2
XFILLER_0_94_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06659_ final_design.cpu.reg_window\[26\] final_design.cpu.reg_window\[58\] net952
+ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout907_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ net465 _04103_ _04257_ _04223_ net456 vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08329_ _03276_ _03277_ _03278_ _03279_ net686 net707 vssd1 vssd1 vccd1 vccd1 _03280_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11340_ net655 net192 vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09024__C1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ net651 _05967_ _05970_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__a21oi_1
X_13010_ net1352 _00241_ net1219 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[30\]
+ sky130_fd_sc_hd__dfrtp_2
X_10222_ final_design.uart.BAUD_counter\[7\] final_design.uart.BAUD_counter\[6\] _05098_
+ final_design.uart.BAUD_counter\[8\] vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_37_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11382__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _05050_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__inv_2
XANTENNA__06484__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input36_A mem_adr_start[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ net1064 final_design.VGA_data_control.v_count\[2\] final_design.VGA_data_control.v_count\[3\]
+ final_design.VGA_data_control.v_count\[1\] vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_54_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09878__A1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 final_design.cpu.reg_window\[10\] vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__dlygate4sd3_1
X_13912_ clknet_leaf_138_clk _01143_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[900\]
+ sky130_fd_sc_hd__dfrtp_1
X_13843_ clknet_leaf_31_clk _01074_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[831\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06458__Y _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11437__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10986_ net1018 _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__nor2_1
X_13774_ clknet_leaf_116_clk _01005_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[762\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14218__1287 vssd1 vssd1 vccd1 vccd1 _14218__1287/HI net1287 sky130_fd_sc_hd__conb_1
XANTENNA__11988__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12725_ _06363_ _06365_ _06361_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_100_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_163_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_163_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11380__X _06067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06864__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12656_ _06315_ net1450 net994 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08833__C net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11607_ net229 net581 net639 vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__and3_1
XANTENNA__11540__B net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12587_ net2431 net1011 net997 final_design.data_from_mem\[5\] vssd1 vssd1 vccd1
+ vccd1 _01280_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06616__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11538_ net680 _05848_ _06124_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold408 final_design.cpu.reg_window\[750\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold419 final_design.cpu.reg_window\[842\] vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09945__B _04863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09015__C1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11469_ net209 net2328 net307 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09566__A0 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13208_ clknet_leaf_132_clk _00439_ net1167 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[196\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14188_ net1258 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XANTENNA__06650__A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13182__RESET_B net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13139_ clknet_leaf_33_clk _00370_ net1129 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13111__RESET_B net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07592__A2 _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 final_design.cpu.reg_window\[267\] vssd1 vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 final_design.cpu.reg_window\[122\] vssd1 vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
X_07700_ final_design.cpu.reg_window\[27\] final_design.cpu.reg_window\[59\] net881
+ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__mux2_1
XANTENNA__09680__B _04598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ _03617_ net603 vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__nand2_4
XANTENNA__10900__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11676__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07631_ _02578_ _02579_ _02580_ _02581_ net694 net713 vssd1 vssd1 vccd1 vccd1 _02582_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11715__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ _01489_ net740 net733 net667 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__and4_2
XANTENNA__12625__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09301_ net498 _04111_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__nand2_2
X_06513_ _01461_ _01462_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__nand2_1
XANTENNA__11979__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09679__Y _04598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07493_ _02130_ _02159_ _02443_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_154_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_154_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11731__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09232_ _03325_ _03355_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__nor2_1
X_06444_ final_design.VGA_data_control.v_count\[7\] final_design.VGA_data_control.v_count\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09201__A _03627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06950__S1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11450__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ net556 net459 _04081_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12038__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08114_ _03052_ _03053_ _03064_ net890 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__a22oi_4
XANTENNA__10403__A2 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09094_ net260 _04016_ _04017_ _04013_ net1030 vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08045_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__nor2_2
XANTENNA__10781__S net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold920 final_design.cpu.reg_window\[370\] vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold931 final_design.cpu.reg_window\[320\] vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1132_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold942 final_design.cpu.reg_window\[613\] vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 final_design.cpu.reg_window\[469\] vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08251__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold964 final_design.cpu.reg_window\[777\] vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 final_design.cpu.reg_window\[109\] vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold986 final_design.cpu.reg_window\[593\] vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11178__A net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold997 final_design.cpu.reg_window\[828\] vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09996_ _02738_ _03594_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout1018_X net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07943__X _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ _03885_ _03887_ net258 vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08207__S1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout857_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09590__B _04508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10810__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _03775_ _03825_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11625__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07829_ final_design.cpu.reg_window\[277\] final_design.cpu.reg_window\[309\] net884
+ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout645_X net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ final_design.CPU_instr_adr\[19\] _03903_ net1070 vssd1 vssd1 vccd1 vccd1
+ _05573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10771_ _05403_ _05502_ _05505_ _05506_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__a211o_1
XANTENNA__12092__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_145_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_145_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12510_ _06172_ net349 net328 net1504 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_142_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13490_ clknet_leaf_26_clk _00721_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[478\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09111__A final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12441_ net1931 net218 net335 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08143__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09796__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12372_ net2207 net220 net270 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_157_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14111_ clknet_leaf_53_clk _01308_ net1159 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_11323_ net600 net196 vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__and2_2
XANTENNA__10691__S net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10059__A1_N _04571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14042_ clknet_leaf_49_clk _00034_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11254_ _02030_ net649 _05954_ _05955_ net661 vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08161__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11088__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _05083_ net811 _05091_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_128_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11185_ _05855_ _05894_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10136_ _01383_ final_design.VGA_data_control.state\[1\] _05039_ vssd1 vssd1 vccd1
+ vccd1 final_design.VGA_data_control.next_state\[0\] sky130_fd_sc_hd__a21o_1
XANTENNA__09781__A _04697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10067_ _04198_ _04983_ _04984_ _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__nand4_1
XANTENNA__11658__A1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11122__A3 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09929__C_N _04847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10330__B2 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_5__f_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload1_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13826_ clknet_leaf_20_clk _01057_ net1103 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[814\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09079__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07709__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12083__A1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_136_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_136_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13757_ clknet_leaf_12_clk _00988_ net1094 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[745\]
+ sky130_fd_sc_hd__dfrtp_1
X_10969_ _04385_ net249 net677 vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06837__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12708_ final_design.VGA_data_control.v_count\[3\] _06348_ _06347_ vssd1 vssd1 vccd1
+ vccd1 _06349_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_128_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13688_ clknet_leaf_131_clk _00919_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[676\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07240__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08039__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ final_design.VGA_data_control.ready_data\[7\] net1033 net988 final_design.data_from_mem\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold205 final_design.cpu.reg_window\[731\] vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07747__Y _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold216 final_design.cpu.reg_window\[472\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold227 final_design.cpu.reg_window\[721\] vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__A0 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold238 final_design.cpu.reg_window\[188\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07476__A _02390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold249 net143 vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09850_ net98 _04180_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout707 net716 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_4
Xfanout718 net724 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__clkbuf_8
Xfanout729 _01720_ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _03671_ _03751_ _03672_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__a21boi_1
X_09781_ _04697_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nor2_1
X_06993_ final_design.cpu.reg_window\[271\] final_design.cpu.reg_window\[303\] net910
+ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__mux2_1
X_08732_ _03681_ _03682_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__and2_1
XANTENNA__12321__S net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08663_ _01999_ _02061_ _02029_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10321__B2 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07614_ final_design.cpu.reg_window\[797\] final_design.cpu.reg_window\[829\] net883
+ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__mux2_1
X_08594_ final_design.cpu.reg_window\[576\] final_design.cpu.reg_window\[608\] net871
+ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12074__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07545_ final_design.cpu.reg_window\[735\] final_design.cpu.reg_window\[767\] net927
+ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_127_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout340_A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout438_A _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10624__A2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07476_ _02390_ _02394_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06555__A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06427_ net73 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11180__B net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09215_ _02997_ _03029_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout605_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09146_ net468 _04064_ _04062_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11585__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09077_ net628 _04001_ _03999_ net261 vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_20_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10805__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08028_ final_design.cpu.reg_window\[851\] final_design.cpu.reg_window\[883\] net828
+ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__mux2_1
XANTENNA__10411__A2_N _05188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold750 final_design.cpu.reg_window\[86\] vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout974_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11337__B1 _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 final_design.cpu.reg_window\[412\] vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout595_X net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold772 final_design.cpu.reg_window\[599\] vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
X_14217__1286 vssd1 vssd1 vccd1 vccd1 _14217__1286/HI net1286 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_9_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold783 final_design.cpu.reg_window\[955\] vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 final_design.cpu.reg_window\[689\] vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08753__A1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ _04896_ _04897_ _04890_ _04894_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__a211o_1
XANTENNA__11195__X _05904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ net1332 _00221_ net1161 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07325__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11941_ _06142_ net283 net408 net2271 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11872_ net193 net563 vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__and2_1
X_13611_ clknet_leaf_16_clk _00842_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[599\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10823_ net1066 _05553_ net1013 final_design.CPU_instr_adr\[18\] vssd1 vssd1 vccd1
+ vccd1 _05557_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_49_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_118_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07167__S1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13542_ clknet_leaf_169_clk _00773_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[530\]
+ sky130_fd_sc_hd__dfrtp_1
X_10754_ _01363_ _03930_ net1070 vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__mux2_1
XANTENNA__13803__RESET_B net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07492__A1 _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10685_ _05410_ _05411_ _05408_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_129_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13473_ clknet_leaf_162_clk _00704_ net1107 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[461\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07995__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09769__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12424_ _06111_ net356 net341 net1894 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_97_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08680__A _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12355_ net2462 net362 net355 _06039_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11306_ net651 _05998_ _06001_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__a21o_1
X_12286_ net566 _06216_ net505 net368 net2267 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_147_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08419__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10434__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11237_ net598 _05939_ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__and3_2
X_14025_ clknet_leaf_85_clk _01256_ net1238 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1013\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_112_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12540__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ final_design.reqhand.data_from_UART\[3\] final_design.data_from_mem\[3\]
+ net249 vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10551__A1 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10551__B2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ final_design.VGA_data_control.v_count\[6\] _05026_ vssd1 vssd1 vccd1 vccd1
+ _05029_ sky130_fd_sc_hd__or2_1
XANTENNA__11546__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12141__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06850__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11099_ _05801_ _05805_ _05804_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10450__A _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11265__B net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12056__A1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13809_ clknet_leaf_109_clk _01040_ net1232 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[797\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_109_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07330_ net771 _02280_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07261_ net673 _01598_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_119_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09000_ _02452_ _02454_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__nand2_1
XANTENNA__08107__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12359__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_07192_ final_design.cpu.reg_window\[841\] final_design.cpu.reg_window\[873\] net925
+ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__mux2_1
XANTENNA__11567__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07235__A1 _01568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10625__A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__B net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12316__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09902_ _04340_ _04817_ _04818_ _04277_ _04118_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10912__X _05642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout504 _06264_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout526 net527 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_6
XANTENNA__12531__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout537 _02211_ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__buf_2
X_09833_ _03228_ net442 vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__nor2_1
Xfanout548 _01908_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_2
XANTENNA_fanout290_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11456__A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__S net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _04394_ _04396_ net480 vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__mux2_1
X_06976_ final_design.cpu.reg_window\[976\] final_design.cpu.reg_window\[1008\] net957
+ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__mux2_1
X_08715_ final_design.CPU_instr_adr\[25\] _01660_ vssd1 vssd1 vccd1 vccd1 _03666_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11098__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12295__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09695_ net736 _04613_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__and2_1
XANTENNA__11890__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08646_ net557 _02733_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_7_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08577_ final_design.cpu.reg_window\[384\] final_design.cpu.reg_window\[416\] net862
+ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout722_A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ final_design.cpu.reg_window\[287\] final_design.cpu.reg_window\[319\] net923
+ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13285__RESET_B net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07474__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07459_ final_design.cpu.reg_window\[960\] final_design.cpu.reg_window\[992\] net951
+ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__mux2_1
XANTENNA__11270__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10470_ net36 _05220_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09129_ _02771_ _03594_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_40_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12140_ net215 net2501 net384 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__mux2_1
XANTENNA__09883__X _04802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout977_X net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12071_ net577 _05929_ net512 net393 net2022 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold580 final_design.cpu.reg_window\[1001\] vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 final_design.cpu.reg_window\[85\] vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _05735_ _05746_ net55 vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__o21bai_1
XANTENNA__12522__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10533__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10533__B2 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__B net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ net1323 _00210_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11924_ _06127_ net288 net410 net2425 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06894__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07162__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _06105_ net282 net520 net1864 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__a22o_1
XANTENNA_output105_A net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10806_ _05522_ _05525_ _05540_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__or3_1
XFILLER_0_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11786_ net2387 net413 net285 _05952_ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10429__B _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13525_ clknet_leaf_53_clk _00756_ net1152 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[513\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10737_ net1066 _05471_ net1013 final_design.CPU_instr_adr\[14\] vssd1 vssd1 vccd1
+ vccd1 _05475_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_24_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ clknet_leaf_112_clk _00687_ net1211 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[444\]
+ sky130_fd_sc_hd__dfrtp_1
X_10668_ net69 final_design.VGA_adr\[8\] _05407_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11549__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12407_ _06105_ net348 net339 net1844 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_114_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12210__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12136__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10599_ net65 _05330_ _05342_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_11_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13387_ clknet_leaf_20_clk _00618_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[375\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08965__B2 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12937__RESET_B net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12338_ net2314 net360 net347 _05911_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09953__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12269_ net568 _06199_ net505 net368 net2363 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__a32o_1
X_14008_ clknet_leaf_132_clk _01239_ net1177 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[996\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12513__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09390__A1 _04308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06830_ final_design.cpu.reg_window\[533\] final_design.cpu.reg_window\[565\] net963
+ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12277__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06761_ final_design.cpu.reg_window\[663\] final_design.cpu.reg_window\[695\] net911
+ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__mux2_1
X_08500_ _02330_ net625 vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__nor2_1
X_06692_ net771 _01642_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__or2_1
X_09480_ _04395_ _04398_ net490 vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13725__RESET_B net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08431_ _03378_ _03379_ _03380_ _03381_ net682 net699 vssd1 vssd1 vccd1 vccd1 _03382_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12029__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11723__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06900__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08362_ final_design.cpu.reg_window\[903\] final_design.cpu.reg_window\[935\] net833
+ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14216__1285 vssd1 vssd1 vccd1 vccd1 _14216__1285/HI net1285 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_22_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07313_ _02260_ _02261_ _02262_ _02263_ net774 net796 vssd1 vssd1 vccd1 vccd1 _02264_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07456__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08293_ net726 _03243_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07244_ final_design.cpu.reg_window\[263\] final_design.cpu.reg_window\[295\] net916
+ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08524__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07175_ net895 _02119_ _02125_ _02107_ _02113_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_147_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12046__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout303_A net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12752__A2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11960__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11885__S net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout301 net302 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout312 net314 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_8
Xfanout323 net324 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_8
Xfanout334 _06283_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11712__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 net346 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07916__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11186__A net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout356 net357 vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_4
XANTENNA__09381__A1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ net490 _04459_ _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__a21o_1
Xfanout367 _06275_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1000_X net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout378 net379 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_8
Xfanout389 _06265_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_6
XANTENNA__12268__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ net484 _04664_ _04665_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a21oi_1
X_06959_ _01909_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout937_A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11914__A final_design.cpu.reg_window\[411\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ _04595_ _04596_ _04594_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07603__S net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08341__C1 _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__Y _05901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11633__B net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ net606 _03065_ _03041_ _02059_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11640_ net571 net420 _06177_ net299 net1899 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__a32o_1
XFILLER_0_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11779__B1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_2_0_clk_X clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10046__A3 _04597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11571_ net437 net593 _06141_ net306 net1500 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__a32o_1
XFILLER_0_107_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13310_ clknet_leaf_146_clk _00541_ net1127 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[298\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10451__B1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10522_ net94 final_design.VGA_adr\[2\] vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13241_ clknet_leaf_168_clk _00472_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[229\]
+ sky130_fd_sc_hd__dfrtp_1
X_10453_ net1427 net1047 _05210_ net248 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input66_A mem_adr_start[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ net1 net1045 vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13172_ clknet_4_9__leaf_clk _00403_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[160\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06958__B1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11951__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12123_ net1741 net183 net390 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__mux2_1
XANTENNA__06889__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12054_ net2386 net184 net399 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__mux2_1
X_11005_ _05729_ _05730_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout890 _01687_ vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12956_ clknet_leaf_50_clk _00194_ net1155 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07686__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11907_ net195 net2131 net274 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ clknet_leaf_87_clk _00125_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_56_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ net185 net2192 net269 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__mux2_1
XANTENNA__09427__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07438__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11769_ net230 net2298 net414 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_40_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ clknet_leaf_106_clk _00739_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[496\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13439_ clknet_leaf_136_clk _00670_ net1170 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[427\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08938__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10745__B2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ final_design.CPU_instr_adr\[17\] _03792_ vssd1 vssd1 vccd1 vccd1 _03917_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07931_ final_design.cpu.reg_window\[854\] final_design.cpu.reg_window\[886\] net822
+ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__mux2_1
XANTENNA__12498__A1 _05869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13977__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ final_design.cpu.reg_window\[20\] final_design.cpu.reg_window\[52\] net867
+ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__mux2_1
X_09601_ _02705_ net447 net444 _02703_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__o22a_1
X_06813_ _01760_ _01761_ _01762_ _01763_ net789 net794 vssd1 vssd1 vccd1 vccd1 _01764_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_127_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07793_ _02740_ _02741_ _02742_ _02743_ net692 net714 vssd1 vssd1 vccd1 vccd1 _02744_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09115__A1 final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09532_ _04429_ _04450_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__and2_1
X_06744_ final_design.cpu.reg_window\[471\] final_design.cpu.reg_window\[503\] net934
+ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__mux2_1
XANTENNA__08519__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08746__C _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ _02735_ _04281_ _02769_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__a21oi_1
X_06675_ net898 _01619_ _01625_ _01612_ _01613_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__a32oi_1
XANTENNA_fanout253_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08414_ _03361_ _03362_ _03363_ _03364_ net684 net704 vssd1 vssd1 vccd1 vccd1 _03365_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09394_ net496 _04312_ _04231_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09418__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08345_ _03103_ _03166_ _03231_ _03295_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__and4_2
XANTENNA_fanout420_A net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1162_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_31_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout518_A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08276_ net616 _03224_ _03225_ net540 vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07227_ final_design.cpu.reg_window\[840\] final_design.cpu.reg_window\[872\] net942
+ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout306_X net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1048_X net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07158_ final_design.cpu.reg_window\[10\] final_design.cpu.reg_window\[42\] net935
+ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux2_1
XANTENNA__11933__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07089_ final_design.cpu.reg_window\[12\] final_design.cpu.reg_window\[44\] net927
+ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__mux2_1
XANTENNA__11187__Y _05897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1107 net1111 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_2
Xfanout1118 net1128 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1129 net1130 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_98_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09354__A1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout186 _06052_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_2
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_2
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12810_ net1364 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_87_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13790_ clknet_leaf_146_clk _01021_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[778\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12741_ final_design.VGA_adr\[3\] net808 _06380_ net967 vssd1 vssd1 vccd1 vccd1 _01350_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12661__B2 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06457__B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10672__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12672_ _06323_ net1410 net991 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11623_ net217 net639 vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__and2_1
XANTENNA__11216__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08672__B _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11554_ net219 net642 vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__and2_1
XANTENNA__09290__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10505_ _05251_ _05253_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_150_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ net189 net2456 net309 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13224_ clknet_leaf_118_clk _00455_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[212\]
+ sky130_fd_sc_hd__dfrtp_1
X_10436_ _03022_ net601 vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__or2_1
XANTENNA_input69_X net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11924__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13155_ clknet_leaf_7_clk _00386_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[143\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10367_ net9 net1036 net1019 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1
+ _00120_ sky130_fd_sc_hd__o22a_1
X_12106_ net2074 net213 net390 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__mux2_1
X_10298_ final_design.VGA_data_control.data_to_VGA\[3\] final_design.VGA_data_control.data_to_VGA\[2\]
+ final_design.VGA_data_control.data_to_VGA\[1\] final_design.VGA_data_control.data_to_VGA\[0\]
+ final_design.VGA_data_control.h_count\[1\] final_design.VGA_data_control.h_count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__mux4_1
X_13086_ clknet_leaf_21_clk _00317_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14215__1284 vssd1 vssd1 vccd1 vccd1 _14215__1284/HI net1284 sky130_fd_sc_hd__conb_1
XANTENNA__10442__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08148__A2 _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12037_ net1515 net215 net396 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09896__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11554__A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13317__RESET_B net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13988_ clknet_leaf_106_clk _01219_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[976\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07243__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11273__B net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ clknet_leaf_67_clk _00177_ net1223 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07470__C _02095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06460_ _01405_ _01412_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_122_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09959__A net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08130_ final_design.cpu.reg_window\[141\] final_design.cpu.reg_window\[173\] net830
+ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12952__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__A0 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08061_ final_design.cpu.reg_window\[786\] final_design.cpu.reg_window\[818\] net818
+ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07012_ final_design.cpu.reg_window\[527\] final_design.cpu.reg_window\[559\] net907
+ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11915__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10055__D _04884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11729__A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12324__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08963_ _03794_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__or2_1
XANTENNA__11448__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06493__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07914_ _01722_ net618 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__nor2_1
X_08894_ _03664_ _03772_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09887__A2 _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12340__B1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07845_ _02790_ _02795_ net723 vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout370_A net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout468_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ final_design.cpu.reg_window\[600\] final_design.cpu.reg_window\[632\] net865
+ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__mux2_1
XANTENNA__06558__A _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09639__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07153__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ net553 net552 net551 net549 net453 net462 vssd1 vssd1 vccd1 vccd1 _04434_
+ sky130_fd_sc_hd__mux4_2
X_06727_ final_design.cpu.reg_window\[792\] final_design.cpu.reg_window\[824\] net950
+ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12643__B2 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_X net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout635_A _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07745__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06992__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09446_ net474 _04223_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__or2_1
X_06658_ final_design.cpu.reg_window\[90\] final_design.cpu.reg_window\[122\] net953
+ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout802_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09377_ net455 _04223_ _04293_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06589_ net561 _01538_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08328_ final_design.cpu.reg_window\[904\] final_design.cpu.reg_window\[936\] net838
+ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__mux2_1
XANTENNA__10957__A1 _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09811__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10957__B2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ final_design.cpu.reg_window\[138\] final_design.cpu.reg_window\[170\] net852
+ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__mux2_1
XANTENNA__12159__A0 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09621__A_N _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11270_ _01967_ net649 _05968_ _05969_ net661 vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__A0 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11198__X _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ net2550 _05099_ _05101_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06740__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11382__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07328__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10152_ _01384_ _05048_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06484__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10083_ final_design.VGA_data_control.v_count\[8\] _04998_ _01404_ vssd1 vssd1 vccd1
+ vccd1 _04999_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_54_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 final_design.cpu.reg_window\[3\] vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08535__C1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13911_ clknet_leaf_137_clk _01142_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[899\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08667__B _02061_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13410__RESET_B net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ clknet_leaf_39_clk _01073_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[830\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13773_ clknet_leaf_139_clk _01004_ net1179 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[761\]
+ sky130_fd_sc_hd__dfrtp_1
X_10985_ _05690_ _05709_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12724_ final_design.VGA_data_control.v_count\[1\] _06364_ vssd1 vssd1 vccd1 vccd1
+ _06365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ final_design.VGA_data_control.ready_data\[15\] net1035 net990 final_design.data_from_mem\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12398__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11606_ net228 net639 vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__and2_1
XFILLER_0_170_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12586_ net2575 net1011 net997 final_design.data_from_mem\[4\] vssd1 vssd1 vccd1
+ vccd1 _01279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11537_ net815 _02359_ net817 vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__or3b_1
XFILLER_0_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold409 final_design.cpu.reg_window\[493\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
X_11468_ net210 net646 vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_78_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13207_ clknet_leaf_144_clk _00438_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[195\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09566__A1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ _03224_ _05190_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__nor2_4
X_14187_ net133 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12144__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ net669 _03781_ net746 vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07238__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ clknet_leaf_44_clk _00369_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13069_ clknet_leaf_127_clk _00300_ net1192 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[57\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1109 final_design.cpu.reg_window\[824\] vssd1 vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08858__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11676__A2 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10900__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11284__A _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07630_ final_design.cpu.reg_window\[412\] final_design.cpu.reg_window\[444\] net875
+ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__mux2_1
X_07561_ net752 _01481_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12625__B2 final_design.data_from_mem\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09300_ net497 _04112_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__nor2_2
X_06512_ _01461_ _01462_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07492_ _02155_ _02157_ _02439_ _02440_ _02187_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__o221a_1
XFILLER_0_91_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09231_ _03388_ _03421_ _03389_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06443_ final_design.vga.v_current_state\[1\] final_design.vga.v_current_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__and2b_1
XANTENNA__11731__B net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12319__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09162_ net623 _03550_ _01658_ _02423_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__a211o_1
XANTENNA__09201__B _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10347__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08113_ _03058_ _03063_ net719 vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__mux2_1
XANTENNA__07002__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ net629 _04014_ net260 vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08044_ net617 _02991_ _02992_ net551 vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__a211oi_4
Xhold910 final_design.cpu.reg_window\[877\] vssd1 vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 final_design.cpu.reg_window\[272\] vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold932 final_design.cpu.reg_window\[269\] vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 final_design.cpu.reg_window\[1012\] vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 final_design.cpu.reg_window\[224\] vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12054__S net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1125_A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 final_design.cpu.reg_window\[147\] vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 final_design.cpu.reg_window\[647\] vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 final_design.cpu.reg_window\[949\] vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 final_design.cpu.reg_window\[126\] vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ net321 _04684_ _04781_ net319 _04913_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout585_A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11893__S net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _03886_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__inv_2
XANTENNA__09871__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _03659_ _03774_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout752_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11194__A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07828_ final_design.cpu.reg_window\[341\] final_design.cpu.reg_window\[373\] net884
+ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07759_ final_design.cpu.reg_window\[472\] final_design.cpu.reg_window\[504\] net868
+ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10770_ _05440_ _05501_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12296__Y _06275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_143_Left_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07611__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11641__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09429_ _04225_ _04343_ _04339_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__o21a_1
XANTENNA__14027__RESET_B net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14214__1283 vssd1 vssd1 vccd1 vccd1 _14214__1283/HI net1283 sky130_fd_sc_hd__conb_1
X_12440_ net1764 net220 net335 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__mux2_1
XANTENNA__09886__X _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08143__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12371_ net1824 net245 net270 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14110_ clknet_leaf_52_clk _01307_ net1151 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.data_from_UART\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_11322_ _04597_ _06015_ net659 vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__mux2_4
XFILLER_0_105_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14229__1294 vssd1 vssd1 vccd1 vccd1 _14229__1294/HI net1294 sky130_fd_sc_hd__conb_1
X_14041_ clknet_leaf_51_clk _00033_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11253_ net744 _03950_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_56_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_152_Left_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12552__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ final_design.uart.BAUD_counter\[1\] final_design.uart.BAUD_counter\[0\] vssd1
+ vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_128_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11184_ final_design.reqhand.data_from_UART\[5\] final_design.data_from_mem\[5\]
+ net249 vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10135_ final_design.VGA_data_control.state\[1\] _01402_ _05038_ final_design.VGA_data_control.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__and4b_1
XANTENNA__08678__A _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07582__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ _04550_ _04551_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__nand2_1
XANTENNA__11658__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13825_ clknet_leaf_154_clk _01056_ net1116 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[813\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12607__B2 final_design.data_from_mem\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08684__Y _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_161_Left_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07709__S1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13756_ clknet_leaf_152_clk _00987_ net1117 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[744\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10968_ net2556 net1041 _05694_ _05695_ vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12707_ _01391_ _06338_ _06343_ _06346_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06837__A2 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11291__B1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13687_ clknet_leaf_137_clk _00918_ net1172 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[675\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10448__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12139__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10899_ _05593_ _05612_ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08039__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12638_ _06306_ net1486 net992 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12795__26 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__inv_2
XFILLER_0_127_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12569_ net2375 _06289_ _06286_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold206 final_design.cpu.reg_window\[712\] vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06661__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__S0 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold217 final_design.cpu.reg_window\[464\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold228 final_design.cpu.reg_window\[688\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_170_Left_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09539__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14239_ net1304 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_169_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07476__B _02394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 final_design.cpu.reg_window\[845\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_169_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12543__B1 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout708 net709 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_4
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout719 net720 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _03675_ _03676_ _03749_ _03673_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_42_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09780_ _04187_ _04698_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06992_ final_design.cpu.reg_window\[335\] final_design.cpu.reg_window\[367\] net910
+ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__mux2_1
X_08731_ final_design.CPU_instr_adr\[14\] _02000_ vssd1 vssd1 vccd1 vccd1 _03682_
+ sky130_fd_sc_hd__or2_1
XANTENNA__06600__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08662_ _01998_ _02029_ _02062_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__or3_2
XANTENNA__07846__A1_N net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07613_ final_design.cpu.reg_window\[861\] final_design.cpu.reg_window\[893\] net880
+ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__mux2_1
X_08593_ final_design.cpu.reg_window\[640\] final_design.cpu.reg_window\[672\] net871
+ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09475__A0 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07544_ net761 _02494_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__or2_1
XANTENNA__08527__S net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__A1 final_design.VGA_data_control.v_count\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09570__S0 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07475_ _02419_ _02424_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12049__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout333_A net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06555__B _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1075_A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ _02803_ _02836_ _04128_ _04132_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_9_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06426_ final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11888__S net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09145_ net532 net459 _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout500_A _06264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_X net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11585__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09076_ final_design.CPU_instr_adr\[6\] _03785_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_20_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08262__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06461__A0 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08027_ net725 _02977_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1030_X net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold740 final_design.cpu.reg_window\[832\] vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11337__A1 _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold751 final_design.cpu.reg_window\[792\] vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1128_X net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold762 final_design.cpu.reg_window\[537\] vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12534__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold773 final_design.cpu.reg_window\[136\] vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 final_design.cpu.reg_window\[398\] vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 final_design.cpu.reg_window\[443\] vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout588_X net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__A2 _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ _03327_ _04895_ _04046_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_51_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13002__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ final_design.CPU_instr_adr\[23\] net1028 _03867_ _03871_ vssd1 vssd1 vccd1
+ vccd1 _00234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08505__A2 _03450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11940_ _06141_ net294 net411 net1976 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11871_ net425 net195 net563 net520 net1895 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13610_ clknet_leaf_1_clk _00841_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[598\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10822_ net977 _05555_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12065__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09466__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10076__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13541_ clknet_leaf_4_clk _00772_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[529\]
+ sky130_fd_sc_hd__dfrtp_1
X_10753_ _05484_ _05488_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13472_ clknet_leaf_35_clk _00703_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[460\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input96_A memory_size[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ net251 _04654_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__and2b_1
XANTENNA__07492__A2 _02157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12423_ _06245_ net503 net341 net2384 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10379__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08680__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08172__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12354_ net2358 net361 net345 _06032_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11305_ _01853_ net649 _05999_ _06000_ net661 vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_75_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12285_ net596 _06215_ net519 net371 net2321 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__a32o_1
XANTENNA__11328__A1 final_design.data_from_mem\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12525__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input51_X net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14024_ clknet_leaf_119_clk _01255_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1012\]
+ sky130_fd_sc_hd__dfrtp_1
X_11236_ _04676_ net661 vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ net740 _04022_ _05878_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_143_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10118_ _05003_ _05027_ _05028_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[5\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__11546__B net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11098_ _04177_ net252 _04990_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06850__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10450__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10049_ _04452_ _04454_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08052__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11265__C net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11562__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ clknet_leaf_110_clk _01039_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[796\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08347__S net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07251__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11264__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13739_ clknet_leaf_17_clk _00970_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[727\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11803__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07260_ _02193_ _02199_ _02210_ net895 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_6_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08107__S1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07191_ net760 _02135_ net755 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11567__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08437__A_N net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10625__B final_design.VGA_adr\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12516__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09901_ _04124_ _04812_ _04813_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout505 net508 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_4
Xfanout516 net517 vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_4
X_09832_ net69 _04182_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__xnor2_1
Xfanout527 _06119_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout538 _02184_ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_2
XANTENNA__12531__A3 _06268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_141_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 _01880_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07426__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213__1282 vssd1 vssd1 vccd1 vccd1 _14213__1282/HI net1282 sky130_fd_sc_hd__conb_1
XANTENNA__11456__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ _03585_ _03589_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__nand2_1
X_06975_ final_design.cpu.reg_window\[784\] final_design.cpu.reg_window\[816\] net957
+ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout283_A _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ final_design.CPU_instr_adr\[25\] _01660_ vssd1 vssd1 vccd1 vccd1 _03665_
+ sky130_fd_sc_hd__nor2_1
X_09694_ net448 _04600_ _04610_ _04612_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__o22a_2
XANTENNA__08499__B2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08645_ _02772_ _03593_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_156_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout548_A _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14228__1293 vssd1 vssd1 vccd1 vccd1 _14228__1293/HI net1293 sky130_fd_sc_hd__conb_1
XFILLER_0_7_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08576_ final_design.cpu.reg_window\[448\] final_design.cpu.reg_window\[480\] net863
+ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__mux2_1
XANTENNA__08257__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10058__A1 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07527_ final_design.cpu.reg_window\[351\] final_design.cpu.reg_window\[383\] net926
+ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout336_X net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout715_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1078_X net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07458_ final_design.cpu.reg_window\[768\] final_design.cpu.reg_window\[800\] net951
+ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06409_ final_design.CPU_instr_adr\[14\] vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07389_ final_design.cpu.reg_window\[194\] final_design.cpu.reg_window\[226\] net939
+ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11411__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09128_ net666 _04045_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__nand2_2
XFILLER_0_162_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09059_ _03787_ _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12507__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12070_ net2376 net392 net500 _05922_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__a22o_1
Xhold570 final_design.cpu.reg_window\[725\] vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold581 final_design.cpu.reg_window\[389\] vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold592 final_design.cpu.reg_window\[847\] vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08499__Y _03450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11021_ net978 _05743_ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__o21a_1
XANTENNA__11647__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__A1 _04109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11730__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07563__C net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12972_ net1322 _00209_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.CPU_instr_adr\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09687__A0 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07860__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11923_ _06126_ net286 net409 net2064 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__a22o_1
XANTENNA__07162__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14042__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09123__Y _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ _06104_ net284 net521 net2138 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07071__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10805_ net44 _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11785_ net2546 net414 _06232_ net432 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11797__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13524_ clknet_leaf_103_clk _00755_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[512\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10736_ net977 _05473_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_24_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input99_X net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13455_ clknet_leaf_92_clk _00686_ net1234 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[443\]
+ sky130_fd_sc_hd__dfrtp_1
X_10667_ net69 final_design.VGA_adr\[8\] _05407_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11549__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12406_ _06104_ net351 net340 net2066 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13386_ clknet_leaf_3_clk _00617_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[374\]
+ sky130_fd_sc_hd__dfrtp_1
X_10598_ _05330_ _05342_ net65 vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_114_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07100__A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__clkbuf_4
XANTENNA__07622__C1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12337_ net2280 net361 net347 _05905_ vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12268_ net584 _06198_ net514 net370 net2015 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14007_ clknet_leaf_143_clk _01238_ net1189 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[995\]
+ sky130_fd_sc_hd__dfrtp_1
X_11219_ final_design.data_from_mem\[9\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1 _05925_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_162_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12152__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ net586 _06127_ net515 net378 net1882 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__a32o_1
XANTENNA__07246__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11991__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11844__X _06239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06760_ final_design.cpu.reg_window\[727\] final_design.cpu.reg_window\[759\] net911
+ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__mux2_1
XANTENNA__11485__A0 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06691_ _01638_ _01639_ _01640_ _01641_ net786 net804 vssd1 vssd1 vccd1 vccd1 _01642_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11292__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08430_ final_design.cpu.reg_window\[517\] final_design.cpu.reg_window\[549\] net821
+ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06900__A1 _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ final_design.cpu.reg_window\[967\] final_design.cpu.reg_window\[999\] net832
+ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08102__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07312_ final_design.cpu.reg_window\[645\] final_design.cpu.reg_window\[677\] net904
+ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__mux2_1
XANTENNA__09697__A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08292_ _03239_ _03240_ _03241_ _03242_ net688 net709 vssd1 vssd1 vccd1 vccd1 _03243_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07243_ final_design.cpu.reg_window\[327\] final_design.cpu.reg_window\[359\] net916
+ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12327__S net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07839__S0 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07174_ net768 _02124_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12201__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1038_A _05168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08540__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 _06159_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_4
XANTENNA_fanout498_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7__f_clk_X clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12062__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_8
Xfanout324 net326 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11712__A1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout335 net336 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1205_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout346 net352 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_2
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ net483 _04733_ _04112_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a21o_1
Xfanout357 _06277_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_2
XANTENNA__09381__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 net369 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_8
Xfanout379 _06271_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_4
XANTENNA_fanout665_A _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ net493 _04559_ _04341_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__a21o_1
X_06958_ net792 net671 _01821_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_119_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11914__B _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09677_ _02803_ _02834_ _04330_ net449 vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__a31o_1
XANTENNA__07144__A1 final_design.data_from_mem\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout832_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06889_ final_design.cpu.reg_window\[979\] final_design.cpu.reg_window\[1011\] net908
+ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08628_ net544 _03072_ _03097_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__and3b_1
XFILLER_0_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ final_design.cpu.reg_window\[513\] final_design.cpu.reg_window\[545\] net851
+ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11930__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11570_ net222 net645 vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10521_ _04847_ net252 vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10451__B2 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11141__S net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13240_ clknet_leaf_132_clk _00471_ net1167 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[228\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10452_ _02698_ net602 vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11844__C_N net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13171_ clknet_leaf_34_clk _00402_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[159\]
+ sky130_fd_sc_hd__dfrtp_1
X_10383_ _01372_ _04995_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06958__A1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12122_ net1855 net184 net391 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__mux2_1
XANTENNA_input59_A mem_adr_start[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12053_ net1665 net186 net398 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07066__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ net54 _05728_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout880 net883 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_4
Xfanout891 net892 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__buf_6
Xclkbuf_3_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__08686__A _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07590__A _02504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12955_ clknet_leaf_50_clk _00193_ net1154 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06569__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ net196 net2163 net276 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12886_ clknet_leaf_86_clk _00124_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07686__A2 _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ net187 net2168 net268 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07589__X _02540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ net681 _05850_ _06118_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_155_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10719_ _05438_ _05441_ _05457_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__nand3_1
XFILLER_0_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13507_ clknet_leaf_6_clk _00738_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[495\]
+ sky130_fd_sc_hd__dfrtp_1
X_14212__1281 vssd1 vssd1 vccd1 vccd1 _14212__1281/HI net1281 sky130_fd_sc_hd__conb_1
XANTENNA__12147__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10456__A _02602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11699_ _05965_ net635 vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13438_ clknet_leaf_21_clk _00669_ net1127 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[426\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13369_ clknet_leaf_164_clk _00600_ net1085 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[357\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08360__S net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14227__1292 vssd1 vssd1 vccd1 vccd1 _14227__1292/HI net1292 sky130_fd_sc_hd__conb_1
XFILLER_0_48_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ net725 _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__nor2_1
XANTENNA__12498__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ final_design.cpu.reg_window\[84\] final_design.cpu.reg_window\[116\] net868
+ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__mux2_1
XANTENNA__07374__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09600_ net474 _04211_ _04518_ _04109_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__a211o_1
X_06812_ final_design.cpu.reg_window\[21\] final_design.cpu.reg_window\[53\] net963
+ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07792_ final_design.cpu.reg_window\[409\] final_design.cpu.reg_window\[441\] net863
+ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09531_ net322 _04430_ _04431_ _04449_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__o31ai_2
X_06743_ final_design.cpu.reg_window\[279\] final_design.cpu.reg_window\[311\] net934
+ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09979__X _04898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ _04048_ _04360_ _04361_ _04380_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__a31o_1
X_06674_ net771 _01624_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06547__C net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08413_ final_design.cpu.reg_window\[389\] final_design.cpu.reg_window\[421\] net823
+ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09393_ _04227_ _04295_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_164_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout246_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09418__A3 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08344_ _03259_ _03260_ _03290_ _03292_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__o22a_1
XANTENNA__12422__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12057__S net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11630__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08275_ net604 _03224_ _03200_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__o21a_1
XANTENNA__10433__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout413_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1155_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07226_ net768 _02176_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__or2_1
XFILLER_0_171_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11896__S net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__A2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09051__A1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07157_ final_design.cpu.reg_window\[74\] final_design.cpu.reg_window\[106\] net934
+ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__mux2_1
XANTENNA__08485__S0 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08270__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07088_ final_design.cpu.reg_window\[76\] final_design.cpu.reg_window\[108\] net927
+ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__mux2_1
XANTENNA__11909__B _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1110 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1110_X net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12489__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1119 net1128 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_1__f_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__09354__A2 _04231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 net177 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout187 _06052_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_2
Xfanout198 _06010_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XANTENNA__11449__A0 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07614__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09729_ _03071_ net446 net439 _03068_ _04640_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06738__B net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ _06366_ _06377_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_26_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ final_design.VGA_data_control.ready_data\[23\] net1033 net988 final_design.data_from_mem\[23\]
+ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06971__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11622_ net575 net421 _06168_ net299 net1448 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__a32o_1
XFILLER_0_77_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12413__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08672__C _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11553_ net2258 net303 _06132_ net421 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10424__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10504_ net93 final_design.VGA_adr\[1\] vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__or2_1
Xwire555 _01717_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11484_ net191 net2377 net309 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12177__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13223_ clknet_leaf_8_clk _00454_ net1088 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[211\]
+ sky130_fd_sc_hd__dfrtp_1
X_10435_ net1456 net1040 _05201_ net247 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11924__A1 _06127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13154_ clknet_leaf_29_clk _00385_ net1138 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[142\]
+ sky130_fd_sc_hd__dfrtp_1
X_10366_ net8 net1036 net1019 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1
+ _00119_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_59_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12105_ net1763 net215 net388 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__mux2_1
X_13085_ clknet_leaf_10_clk _00316_ net1091 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[73\]
+ sky130_fd_sc_hd__dfrtp_1
X_10297_ final_design.VGA_data_control.data_to_VGA\[4\] _05013_ _05150_ final_design.VGA_data_control.h_count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a211o_1
XANTENNA__11137__C1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12036_ net1663 net217 net397 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__mux2_1
XANTENNA__11688__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09896__A3 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09305__A _02503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11554__B net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12101__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13987_ clknet_leaf_6_clk _01218_ net1089 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[975\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08305__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09502__C1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12938_ clknet_leaf_68_clk _00176_ net1221 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_157_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11860__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12869_ clknet_leaf_72_clk _00107_ net1244 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12404__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06619__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07816__C1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11612__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__A1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08060_ final_design.cpu.reg_window\[850\] final_design.cpu.reg_window\[882\] net821
+ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12168__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07011_ final_design.cpu.reg_window\[591\] final_design.cpu.reg_window\[623\] net907
+ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__mux2_1
XANTENNA__12992__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10914__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11915__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06603__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11729__B net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09584__A2 _04153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08962_ final_design.CPU_instr_adr\[18\] _03793_ final_design.CPU_instr_adr\[19\]
+ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07913_ net607 _02863_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08893_ _01631_ _01632_ _01662_ _02470_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout196_A _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__A2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07844_ _02791_ _02792_ _02793_ _02794_ net697 net703 vssd1 vssd1 vccd1 vccd1 _02795_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10351__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06839__A _01785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11464__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ final_design.cpu.reg_window\[664\] final_design.cpu.reg_window\[696\] net865
+ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_56_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09514_ _03029_ net446 net442 _03027_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__o221a_1
X_06726_ final_design.cpu.reg_window\[856\] final_design.cpu.reg_window\[888\] net950
+ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09502__X _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09445_ _04362_ _04363_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__nor2_1
XANTENNA__10654__B2 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11851__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06657_ final_design.cpu.reg_window\[154\] final_design.cpu.reg_window\[186\] net952
+ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__mux2_1
XANTENNA__09869__B _04787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout530_A _02502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout628_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08265__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09376_ net493 _04225_ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__or3b_1
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06588_ net752 _01537_ net672 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08327_ final_design.cpu.reg_window\[968\] final_design.cpu.reg_window\[1000\] net839
+ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1060_X net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ final_design.cpu.reg_window\[202\] final_design.cpu.reg_window\[234\] net852
+ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout997_A _06296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07209_ final_design.cpu.reg_window\[328\] final_design.cpu.reg_window\[360\] net921
+ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_65_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09024__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08189_ _03136_ _03137_ _03138_ _03139_ net690 net710 vssd1 vssd1 vccd1 vccd1 _03140_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_160_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10220_ final_design.uart.BAUD_counter\[7\] _05099_ net812 vssd1 vssd1 vccd1 vccd1
+ _05101_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07609__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11639__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11382__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ _05046_ _05048_ _05049_ vssd1 vssd1 vccd1 vccd1 final_design.vga.h_next_count\[2\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_37_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10082_ final_design.VGA_data_control.v_count\[7\] final_design.VGA_data_control.v_count\[5\]
+ final_design.VGA_data_control.v_count\[6\] vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_54_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout952_X net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11655__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13910_ clknet_leaf_124_clk _01141_ net1191 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[898\]
+ sky130_fd_sc_hd__dfrtp_1
X_14211__1280 vssd1 vssd1 vccd1 vccd1 _14211__1280/HI net1280 sky130_fd_sc_hd__conb_1
XFILLER_0_96_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13841_ clknet_leaf_109_clk _01072_ net1232 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[829\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10886__A2_N _05615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13772_ clknet_leaf_125_clk _01003_ net1196 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[760\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ _05694_ _05709_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__or2_1
XANTENNA__10645__A1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11842__A0 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12723_ final_design.VGA_data_control.v_count\[2\] _06359_ vssd1 vssd1 vccd1 vccd1
+ _06364_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_100_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14226__1291 vssd1 vssd1 vccd1 vccd1 _14226__1291/HI net1291 sky130_fd_sc_hd__conb_1
XFILLER_0_155_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12654_ _06314_ net1393 net994 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__mux2_1
XANTENNA__08175__S net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ net230 net2079 net301 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12585_ net1682 net1011 net997 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1
+ vccd1 _01278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11536_ net815 _02358_ net817 vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__and3b_4
XFILLER_0_151_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06771__X _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08471__C1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14255_ net1320 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XANTENNA__09015__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11467_ net211 net2237 net308 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06931__B _01881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ clknet_leaf_129_clk _00437_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[194\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09566__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10418_ net1440 net1043 _05192_ net246 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__a22o_1
X_14186_ net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_1
X_11398_ net428 net580 _06082_ net316 net1639 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07121__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13137_ clknet_leaf_109_clk _00368_ net1230 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[125\]
+ sky130_fd_sc_hd__dfrtp_1
X_10349_ wb_manage.BUSY_O wb_manage.prev_BUSY_O net1037 vssd1 vssd1 vccd1 vccd1 _05170_
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13068_ clknet_leaf_123_clk _00299_ net1191 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12322__A1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ _06221_ net293 net403 net2179 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__a22o_1
XANTENNA__12160__S net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07254__S net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13538__RESET_B net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07560_ _01477_ _01480_ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__nor2_1
XANTENNA__12086__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06511_ final_design.data_from_mem\[6\] net1051 net1007 net1004 vssd1 vssd1 vccd1
+ vccd1 _01462_ sky130_fd_sc_hd__or4_1
XANTENNA__11833__A0 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07491_ _02439_ _02440_ _02187_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__o21a_1
XANTENNA__12396__A net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11504__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09230_ _03423_ _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__nand2_2
X_06442_ final_design.reqhand.current_client\[1\] net1053 _01395_ vssd1 vssd1 vccd1
+ vccd1 _01396_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12389__A1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09161_ _04078_ _04079_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08112_ _03059_ _03060_ _03061_ _03062_ net687 net701 vssd1 vssd1 vccd1 vccd1 _03063_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09092_ _03784_ _04015_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11299__X _05996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08043_ net606 _02991_ _02966_ _01850_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold900 final_design.cpu.reg_window\[621\] vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold911 final_design.cpu.reg_window\[368\] vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout209_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold922 final_design.cpu.reg_window\[273\] vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07429__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12010__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 final_design.cpu.reg_window\[322\] vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 final_design.cpu.reg_window\[388\] vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 final_design.cpu.reg_window\[358\] vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 final_design.cpu.reg_window\[193\] vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 final_design.cpu.reg_window\[68\] vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10021__C1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold988 final_design.cpu.reg_window\[143\] vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ net478 _04411_ _04912_ net320 vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__o211a_1
Xhold999 final_design.cpu.reg_window\[634\] vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1118_A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08945_ final_design.CPU_instr_adr\[21\] _03795_ vssd1 vssd1 vccd1 vccd1 _03886_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__08401__X _03352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ _03823_ _02474_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_32_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07164__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07827_ _02774_ _02775_ _02776_ _02777_ net697 net703 vssd1 vssd1 vccd1 vccd1 _02778_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_84_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout745_A _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ final_design.cpu.reg_window\[280\] final_design.cpu.reg_window\[312\] net868
+ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__mux2_1
XANTENNA__12077__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06709_ net752 _01659_ net672 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__a21o_2
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11824__A0 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07689_ _02637_ _02639_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout912_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12092__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11414__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09428_ _04334_ _04335_ _04346_ net263 vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09359_ net491 _04277_ _04276_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12370_ net1631 net237 net271 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__mux2_1
XANTENNA__09796__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11321_ _01788_ net650 _06014_ net651 _06013_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__a221o_1
XANTENNA__07847__B net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ clknet_leaf_51_clk _00032_ net1155 vssd1 vssd1 vccd1 vccd1 final_design.uart.BAUD_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07339__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ net667 _03944_ net739 vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12001__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10203_ final_design.uart.BAUD_counter\[0\] net811 vssd1 vssd1 vccd1 vccd1 _00006_
+ sky130_fd_sc_hd__and2b_1
X_11183_ net748 _04009_ _05892_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_128_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input41_A mem_adr_start[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ final_design.VGA_data_control.h_count\[0\] _05037_ vssd1 vssd1 vccd1 vccd1
+ _05038_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_73_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08678__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09705__C1 _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ _04510_ _04511_ _04550_ _04551_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_145_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09126__Y _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07074__S net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10866__A1 final_design.CPU_instr_adr\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10866__B2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13824_ clknet_leaf_38_clk _01055_ net1136 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[812\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12068__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07802__S net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10967_ _05673_ _05692_ net1016 vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__o21a_1
X_13755_ clknet_leaf_155_clk _00986_ net1115 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[743\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12083__A3 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12706_ _06340_ _06346_ _06345_ net1064 vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09302__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10898_ _05590_ _05612_ _05611_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__a21bo_1
X_13686_ clknet_leaf_124_clk _00917_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[674\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10448__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12637_ final_design.VGA_data_control.ready_data\[6\] net1033 net988 final_design.data_from_mem\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12568_ final_design.uart.receiving final_design.uart.working_data\[4\] vssd1 vssd1
+ vccd1 vccd1 _06289_ sky130_fd_sc_hd__and2_1
XANTENNA__12240__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11519_ net2151 _06120_ _06121_ net437 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_117_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12155__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10464__A _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12499_ _06160_ net350 net328 net2162 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold207 final_design.cpu.reg_window\[173\] vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07893__S1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold218 final_design.VGA_data_control.ready_data\[23\] vssd1 vssd1 vccd1 vccd1 net1571
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 final_design.cpu.reg_window\[207\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14238_ net1303 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_169_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14169_ clknet_leaf_82_clk _01343_ net1243 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08869__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__buf_4
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06991_ _01940_ _01941_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08730_ final_design.CPU_instr_adr\[14\] _02000_ vssd1 vssd1 vccd1 vccd1 _03681_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08661_ _02545_ _03610_ _02542_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__a21oi_1
X_07612_ _02559_ _02560_ _02561_ _02562_ net696 net715 vssd1 vssd1 vccd1 vccd1 _02563_
+ sky130_fd_sc_hd__mux4_1
X_08592_ final_design.cpu.reg_window\[704\] final_design.cpu.reg_window\[736\] net871
+ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__mux2_1
XANTENNA__06676__X _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06930__C1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07543_ _02490_ _02491_ _02492_ _02493_ net779 net800 vssd1 vssd1 vccd1 vccd1 _02494_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_147_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09475__A1 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12074__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07474_ net749 _01497_ _02420_ _02421_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09213_ _02866_ _04129_ _04130_ _04128_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07581__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06425_ final_design.reqhand.instruction\[20\] vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1068_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ net614 _03549_ _02325_ _02422_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__o211a_1
XANTENNA__12231__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11585__A2 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09075_ _03723_ _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1235_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08026_ _02973_ _02974_ _02975_ _02976_ net683 net704 vssd1 vssd1 vccd1 vccd1 _02977_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold730 final_design.cpu.reg_window\[673\] vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold741 final_design.cpu.reg_window\[654\] vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11337__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout695_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 final_design.cpu.reg_window\[1006\] vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 final_design.cpu.reg_window\[491\] vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09935__C1 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold774 final_design.uart.working_data\[4\] vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1023_X net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold785 final_design.cpu.reg_window\[361\] vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 final_design.cpu.reg_window\[917\] vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07410__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout862_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ _03327_ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ net258 _03869_ net1028 vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10841__A1_N net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08859_ net633 _03806_ _03808_ net261 vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13042__RESET_B net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08910__B1 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11870_ _06017_ net648 net292 net523 net1719 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__a32o_1
XANTENNA__06586__X _01537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10821_ net973 _05553_ _05554_ _04042_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10549__A final_design.CPU_instr_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11144__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10752_ _05467_ _05470_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_137_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13540_ clknet_leaf_98_clk _00771_ net1218 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[528\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12470__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07883__A_N net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13471_ clknet_leaf_135_clk _00702_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[459\]
+ sky130_fd_sc_hd__dfrtp_1
X_10683_ net1454 net1042 net1015 _05423_ vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12422_ _06110_ net355 net341 net2211 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__a22o_1
XANTENNA__12222__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09769__A2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input89_A memory_size[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08306__X _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07324__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12353_ _06236_ net500 net360 net2421 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06988__C1 _01821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11304_ net743 _03902_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__nand2_1
XANTENNA__07069__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12284_ net587 _06214_ net515 net370 net1648 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_75_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14023_ clknet_leaf_9_clk _01254_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1011\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_147_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11235_ net651 _05936_ _05937_ _05938_ net662 vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_112_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input44_X net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ net670 _04020_ net746 vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__a21o_1
XANTENNA__06701__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ net1064 _05023_ final_design.VGA_data_control.v_count\[5\] vssd1 vssd1 vccd1
+ vccd1 _05028_ sky130_fd_sc_hd__a21o_1
XANTENNA__12289__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ _05798_ _05815_ _05814_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11546__C net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10048_ _04529_ _04530_ _04616_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_160_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08052__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 final_design.uart.working_data\[8\] vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11843__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07532__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13807_ clknet_leaf_90_clk _01038_ net1233 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[795\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11562__B net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11999_ _06201_ net282 net400 net1967 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_11_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11264__A1 _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13738_ clknet_leaf_0_clk _00969_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[726\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11281__C _05979_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14249__1314 vssd1 vssd1 vccd1 vccd1 _14249__1314/HI net1314 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_119_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13669_ clknet_leaf_4_clk _00900_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[657\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07190_ net769 _02140_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__or2_1
XANTENNA__12213__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11567__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09983__A _04898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09900_ _03638_ _04087_ _04094_ _03637_ _04811_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a221o_1
XANTENNA__10922__A net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout506 net508 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13553__RESET_B net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ _04745_ _04747_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__xnor2_1
Xfanout517 _06259_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_2
Xfanout539 _02155_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_2
XANTENNA__07943__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06974_ final_design.cpu.reg_window\[848\] final_design.cpu.reg_window\[880\] net957
+ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__mux2_1
X_09762_ _04426_ _04680_ net448 vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a21o_1
XFILLER_0_174_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08713_ _03662_ _03663_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__and2_1
X_09693_ _03164_ _04498_ _04611_ net666 _04045_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12295__A3 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout276_A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ _03040_ _02772_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08538__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08575_ final_design.cpu.reg_window\[256\] final_design.cpu.reg_window\[288\] net863
+ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout443_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1185_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07526_ _01509_ _02476_ _01508_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11899__S net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07457_ final_design.cpu.reg_window\[832\] final_design.cpu.reg_window\[864\] net951
+ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout708_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06408_ final_design.CPU_instr_adr\[15\] vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12204__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07388_ final_design.cpu.reg_window\[2\] final_design.cpu.reg_window\[34\] net946
+ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09127_ net666 _04045_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__and2_4
XFILLER_0_32_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1238_X net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09058_ final_design.CPU_instr_adr\[8\] _03786_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08009_ _02954_ _02959_ net723 vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__mux2_1
XANTENNA__07684__Y _02635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold560 final_design.cpu.reg_window\[1013\] vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10518__B1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09384__A0 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 final_design.cpu.reg_window\[796\] vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net973 _05742_ _05744_ _04042_ net975 vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a221o_1
Xhold582 final_design.cpu.reg_window\[979\] vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 final_design.cpu.reg_window\[166\] vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11647__B _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__A2 _04398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__D net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ clknet_leaf_73_clk net1354 net1244 vssd1 vssd1 vccd1 vccd1 wb_manage.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10978__S net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09687__A1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12286__A3 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ net230 net2490 net410 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__mux2_1
XANTENNA__12691__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08448__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07352__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__S0 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07205__X _02156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11853_ _06103_ net282 net521 net2007 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10804_ net676 _05527_ _05538_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11784_ net656 net565 net214 vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_99_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11797__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13523_ clknet_leaf_32_clk _00754_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[511\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10735_ net973 _05471_ _05472_ _04042_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14011__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10666_ net70 final_design.VGA_adr\[9\] vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__xnor2_1
X_13454_ clknet_leaf_114_clk _00685_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[442\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11549__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ _06103_ net348 net339 net2106 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__a22o_1
X_13385_ clknet_leaf_88_clk _00616_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[373\]
+ sky130_fd_sc_hd__dfrtp_1
X_10597_ _05340_ _05341_ net975 vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12210__A3 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__clkbuf_4
X_12336_ net2301 net360 net344 _05898_ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12433__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ net585 _06197_ net517 net370 net2059 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08178__B2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ net742 _03981_ _05923_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__o21a_1
X_14006_ clknet_leaf_129_clk _01237_ net1176 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[994\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07527__S net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09308__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__A2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12198_ net582 _06126_ net513 net377 net2083 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_162_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11182__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ net660 _05860_ _05862_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12277__A3 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06690_ final_design.cpu.reg_window\[153\] final_design.cpu.reg_window\[185\] net952
+ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08360_ final_design.cpu.reg_window\[775\] final_design.cpu.reg_window\[807\] net856
+ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08102__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07311_ final_design.cpu.reg_window\[709\] final_design.cpu.reg_window\[741\] net904
+ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__mux2_1
XANTENNA__07536__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09697__B _04613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08291_ final_design.cpu.reg_window\[137\] final_design.cpu.reg_window\[169\] net842
+ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11512__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07242_ net768 _02192_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__or2_1
XANTENNA__08093__S net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06606__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07173_ _02120_ _02121_ _02122_ _02123_ net778 net791 vssd1 vssd1 vccd1 vccd1 _02124_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07839__S1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09602__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11960__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout303 net306 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_8
Xfanout314 _06092_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11173__B1 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout393_A _06263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07916__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 _06282_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_6
Xfanout347 net348 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_4
X_09814_ _04618_ _04732_ net472 vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__mux2_1
XANTENNA__09381__A3 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_4
Xfanout369 net371 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10920__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ _04485_ _04663_ net471 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06957_ net894 _01907_ _01896_ _01895_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__12268__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A _05849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09676_ _02834_ _04330_ _02803_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08268__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06888_ final_design.cpu.reg_window\[787\] final_design.cpu.reg_window\[819\] net911
+ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__mux2_1
XANTENNA__06577__A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08627_ _03572_ _03577_ _03167_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08892__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_X net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12425__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08558_ final_design.cpu.reg_window\[577\] final_design.cpu.reg_window\[609\] net851
+ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__mux2_1
XANTENNA__06864__X _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__C1 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11779__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07509_ _01855_ _02459_ _01856_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__o21a_1
X_08489_ final_design.cpu.reg_window\[771\] final_design.cpu.reg_window\[803\] net863
+ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10827__A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11422__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10520_ _05249_ _05264_ _05263_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_42_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10451_ net255 _05209_ net1047 net151 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_94_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11400__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ clknet_leaf_44_clk _00401_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[158\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10382_ net26 net1036 net1019 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1
+ vccd1 _00135_ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12121_ net1874 net186 net390 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13404__RESET_B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11951__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12052_ net2115 net188 net399 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__mux2_1
XANTENNA__09128__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold390 final_design.cpu.reg_window\[914\] vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net54 _05728_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__and2_1
X_14248__1313 vssd1 vssd1 vccd1 vccd1 _14248__1313/HI net1313 sky130_fd_sc_hd__conb_1
XFILLER_0_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10911__B1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 net876 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_4
Xfanout881 net883 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_4
Xfanout892 net893 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12259__A3 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07590__B net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09134__Y _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ clknet_leaf_55_clk _00192_ net1163 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06487__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1090 final_design.cpu.reg_window\[40\] vssd1 vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07766__S0 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06569__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ net197 net1927 net276 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output110_A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ clknet_leaf_87_clk _00123_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08883__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11219__A1 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09798__A _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ net188 net2222 net268 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12416__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11767_ net177 net2232 net417 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__mux2_1
XANTENNA__08635__A2 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_140_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13506_ clknet_leaf_23_clk _00737_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[494\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06646__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10718_ net40 _05456_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11698_ net427 net573 _06207_ net295 net1597 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__a32o_1
XANTENNA__10456__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13437_ clknet_leaf_32_clk _00668_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[425\]
+ sky130_fd_sc_hd__dfrtp_1
X_10649_ _05368_ _05390_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13368_ clknet_leaf_128_clk _00599_ net1178 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[356\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_155_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11942__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ net1672 net195 net364 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13299_ clknet_leaf_31_clk _00530_ net1131 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[287\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09348__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12498__A3 _06268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ net721 _02810_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10902__B1 _05610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ final_design.cpu.reg_window\[85\] final_design.cpu.reg_window\[117\] net963
+ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__mux2_1
X_07791_ final_design.cpu.reg_window\[473\] final_design.cpu.reg_window\[505\] net863
+ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11507__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06742_ final_design.cpu.reg_window\[343\] final_design.cpu.reg_window\[375\] net934
+ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__mux2_1
X_09530_ net263 _04433_ _04445_ _04448_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__and4_1
XANTENNA__08859__C1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _04231_ _04367_ _04372_ _04379_ net264 vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__o2111ai_2
X_06673_ _01620_ _01621_ _01622_ _01623_ net786 net804 vssd1 vssd1 vccd1 vccd1 _01624_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08874__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08412_ final_design.cpu.reg_window\[453\] final_design.cpu.reg_window\[485\] net822
+ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12407__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09392_ _04056_ _04310_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08343_ _03293_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09284__C1 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__B1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout239_A _05890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11630__A1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13915__RESET_B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08274_ _02128_ net616 vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__nor2_1
XANTENNA__10433__A2 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07834__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07225_ _02172_ _02173_ _02174_ _02175_ net782 net791 vssd1 vssd1 vccd1 vccd1 _02176_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout406_A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07156_ net759 _02106_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__or2_1
XANTENNA__08551__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12581__B net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__B1 _06078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08485__S1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11933__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11478__A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11277__A2_N _05947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07087_ _02034_ _02035_ _02036_ _02037_ net779 net800 vssd1 vssd1 vccd1 vccd1 _02038_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1109 net1110 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout775_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08562__A1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07996__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout177 _06089_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_2
Xfanout188 _06045_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
XANTENNA_fanout942_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ final_design.cpu.reg_window\[464\] final_design.cpu.reg_window\[496\] net878
+ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout563_X net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11417__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ _04643_ _04646_ net490 vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ net477 _04458_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_26_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10672__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12670_ _06322_ net1716 net991 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11621_ net220 net639 vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__and2_1
XANTENNA__06971__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10424__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ net574 net244 net642 vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__and3_1
XANTENNA__08027__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09290__A2 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10503_ net93 final_design.VGA_adr\[1\] vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__nor2_1
X_11483_ net191 net647 vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire545 _01995_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_163_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input71_A memory_size[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13222_ clknet_leaf_171_clk _00453_ net1074 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[210\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07866__A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10434_ _02929_ net601 vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_150_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11924__A2 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10365_ net7 net1038 net1021 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1
+ _00118_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13153_ clknet_leaf_159_clk _00384_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[141\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ net1915 net217 net389 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__mux2_1
X_13084_ clknet_leaf_149_clk _00315_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_10296_ final_design.VGA_data_control.h_count\[1\] final_design.VGA_data_control.h_count\[2\]
+ final_design.VGA_data_control.data_to_VGA\[5\] vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__and3b_1
XANTENNA__11137__B1 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12035_ net1645 net219 net396 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__mux2_1
XANTENNA__11688__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06769__X _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10360__B2 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13986_ clknet_leaf_29_clk _01217_ net1140 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[974\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08305__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07106__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12937_ clknet_leaf_67_clk _00175_ net1223 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_166_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_166_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_157_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12868_ clknet_leaf_72_clk _00106_ net1244 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07540__S net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11570__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11819_ net220 net2175 net266 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12158__S net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08164__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11612__A1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09281__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07010_ final_design.cpu.reg_window\[655\] final_design.cpu.reg_window\[687\] net907
+ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__mux2_1
XANTENNA__06680__A _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10914__B _05642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07044__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11915__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08961_ net627 _03896_ net256 vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07912_ _02850_ _02851_ _02862_ net889 vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__a22oi_4
X_08892_ final_design.CPU_instr_adr\[27\] net1029 _03836_ _03838_ vssd1 vssd1 vccd1
+ vccd1 _00238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire531_X net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12340__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07843_ final_design.cpu.reg_window\[533\] final_design.cpu.reg_window\[565\] net884
+ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__mux2_1
XANTENNA__10351__B2 final_design.data_from_mem\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07752__C1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_A _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ final_design.cpu.reg_window\[728\] final_design.cpu.reg_window\[760\] net869
+ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09513_ _03025_ net441 vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__nand2_1
X_06725_ final_design.cpu.reg_window\[920\] final_design.cpu.reg_window\[952\] net950
+ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__mux2_1
XANTENNA__10103__A1 final_design.VGA_data_control.v_count\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_157_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_157_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout356_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06656_ final_design.cpu.reg_window\[218\] final_design.cpu.reg_window\[250\] net953
+ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__mux2_1
X_09444_ net469 _04078_ _04102_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07450__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06587_ net752 _01537_ net672 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ _03485_ _04293_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout523_A _06239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ final_design.cpu.reg_window\[776\] final_design.cpu.reg_window\[808\] net861
+ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14247__1312 vssd1 vssd1 vccd1 vccd1 _14247__1312/HI net1312 sky130_fd_sc_hd__conb_1
XANTENNA__10096__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08257_ final_design.cpu.reg_window\[10\] final_design.cpu.reg_window\[42\] net853
+ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__mux2_1
XANTENNA__09009__C1 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07208_ _02155_ _02157_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06590__A _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08188_ final_design.cpu.reg_window\[398\] final_design.cpu.reg_window\[430\] net852
+ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout892_A net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07139_ _02084_ _02089_ net764 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ final_design.VGA_data_control.h_count\[0\] final_design.VGA_data_control.h_count\[1\]
+ net1062 vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ _01400_ _04996_ _01391_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__and3b_1
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772__3 clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09406__A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11655__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout945_X net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__S net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10342__B2 final_design.data_from_mem\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ clknet_leaf_112_clk _01071_ net1216 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[828\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_148_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_148_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13771_ clknet_leaf_17_clk _01002_ net1099 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[759\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10983_ _05690_ _05694_ _05709_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__nand3_1
XFILLER_0_168_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08394__S0 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11671__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12722_ _06354_ _06362_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06765__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ final_design.VGA_data_control.ready_data\[14\] net1035 net990 final_design.data_from_mem\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__a22o_1
XANTENNA__10287__A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12398__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11604_ net679 _05848_ _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__or3_1
X_12584_ net2476 net1011 net997 final_design.data_from_mem\[2\] vssd1 vssd1 vccd1
+ vccd1 _01277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11535_ net2063 net176 net525 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input74_X net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14254_ net1319 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_150_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08191__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08615__A_N net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11466_ net213 net2488 net309 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__mux2_1
XANTENNA__11358__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13205_ clknet_leaf_40_clk _00436_ net1143 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[193\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10417_ _03257_ _05190_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__nor2_1
X_14185_ clknet_leaf_75_clk final_design.VGA_data_control.next_state\[1\] net1245
+ vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.state\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09566__A3 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11397_ net655 net178 vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__and2_1
XANTENNA__07121__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ clknet_leaf_108_clk _00367_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[124\]
+ sky130_fd_sc_hd__dfrtp_1
X_10348_ wb_manage.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08698__Y _03649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08765__A_N final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__C1 _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10279_ final_design.uart.BAUD_counter\[29\] final_design.uart.BAUD_counter\[28\]
+ _05134_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__and3_1
XANTENNA__12441__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13067_ clknet_leaf_15_clk _00298_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09723__A0 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07535__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ _06220_ net291 net402 net2055 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10333__B2 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07107__Y _02058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12086__A1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_139_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_139_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13969_ clknet_leaf_109_clk _01200_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[957\]
+ sky130_fd_sc_hd__dfrtp_1
X_06510_ net1053 net1006 net1003 final_design.reqhand.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 _01461_ sky130_fd_sc_hd__a31o_1
X_07490_ _02439_ _02440_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_17_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10909__B net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06441_ wb_manage.BUSY_O final_design.reqhand.current_client\[0\] net34 vssd1 vssd1
+ vccd1 vccd1 _01395_ sky130_fd_sc_hd__or3b_2
XFILLER_0_146_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09160_ net623 _03549_ _03523_ _01627_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__a211o_1
XFILLER_0_174_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08111_ final_design.cpu.reg_window\[524\] final_design.cpu.reg_window\[556\] net847
+ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__mux2_1
XANTENNA__11597__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09091_ final_design.CPU_instr_adr\[3\] net1031 final_design.CPU_instr_adr\[4\] vssd1
+ vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11520__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08042_ net606 _02991_ _02966_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_153_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11349__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold901 final_design.cpu.reg_window\[33\] vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 final_design.cpu.reg_window\[704\] vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold923 final_design.cpu.reg_window\[442\] vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 final_design.cpu.reg_window\[314\] vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold945 final_design.cpu.reg_window\[288\] vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 final_design.cpu.reg_window\[630\] vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold967 final_design.cpu.reg_window\[257\] vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 final_design.cpu.reg_window\[459\] vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 final_design.cpu.reg_window\[544\] vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ net471 _04401_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08944_ _03882_ _03884_ net631 vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07953__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1013_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07445__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11475__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _01571_ _01601_ _02473_ net628 vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__a31o_1
XANTENNA__10324__B2 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_A _03485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07826_ final_design.cpu.reg_window\[21\] final_design.cpu.reg_window\[53\] net884
+ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ final_design.cpu.reg_window\[344\] final_design.cpu.reg_window\[376\] net868
+ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout640_A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06708_ final_design.reqhand.instruction\[25\] final_design.data_from_mem\[25\] net985
+ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__mux2_2
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07688_ net613 _02635_ _02611_ net562 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09427_ _02900_ net446 _04344_ _04345_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06639_ final_design.cpu.reg_window\[731\] final_design.cpu.reg_window\[763\] net960
+ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09358_ net478 _04065_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08309_ net619 _03257_ _03258_ net539 vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a211oi_1
X_09289_ _01566_ net560 net459 vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11430__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11320_ final_design.data_from_mem\[21\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06014_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__A2_N net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ final_design.data_from_mem\[13\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1
+ _05953_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10202_ final_design.uart.BAUD_counter_state _05078_ vssd1 vssd1 vccd1 vccd1 _05090_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12552__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11182_ net668 _04006_ net740 vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10133_ final_design.VGA_data_control.h_count\[3\] net1061 final_design.VGA_data_control.h_count\[5\]
+ _05013_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_73_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06862__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07355__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _04962_ _04963_ _04980_ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_145_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10315__B2 final_design.data_from_mem\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10866__A2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09423__X _04342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12068__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ clknet_leaf_137_clk _01054_ net1171 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[811\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12497__A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08694__B _03296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11605__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13754_ clknet_leaf_160_clk _00985_ net1105 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[742\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08186__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10966_ _05673_ _05692_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__nand2_1
XANTENNA__07090__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ net1064 _06344_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__or2_1
XANTENNA__13600__RESET_B net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13685_ clknet_leaf_25_clk _00916_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[673\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11291__A2 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10897_ _04356_ net254 vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12636_ _06305_ net1447 net994 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11579__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12240__A1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ net1406 _06288_ _06286_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__mux2_1
XANTENNA__12436__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11518_ net595 net222 _06116_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__and3_1
XANTENNA__10540__A_N net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10464__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12498_ _05869_ net640 _06268_ net330 net1452 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_117_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold208 final_design.cpu.reg_window\[460\] vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold219 final_design.cpu.reg_window\[186\] vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ net1302 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
X_11449_ net241 net2538 net309 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__mux2_1
XANTENNA__09539__A3 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08747__A1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12543__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14168_ clknet_leaf_79_clk _01342_ net1251 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10554__A1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11751__A0 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10554__B2 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11576__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13119_ clknet_leaf_133_clk _00350_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_84_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12024__X _06259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12171__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14099_ clknet_leaf_83_clk _01296_ net1242 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_06990_ net547 _01939_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__nand2_1
X_14246__1311 vssd1 vssd1 vccd1 vccd1 _14246__1311/HI net1311 sky130_fd_sc_hd__conb_1
XANTENNA__13759__RESET_B net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ _02542_ _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__and2b_1
XANTENNA__06957__X _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ final_design.cpu.reg_window\[669\] final_design.cpu.reg_window\[701\] net878
+ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08591_ net722 _03541_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__or2_1
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11515__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07542_ final_design.cpu.reg_window\[927\] final_design.cpu.reg_window\[959\] net927
+ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08096__S net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06609__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09475__A2 net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07473_ net749 _01497_ _02420_ _02421_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_93_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08683__B1 _02510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09212_ _04130_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10490__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06424_ final_design.data_from_mem\[5\] vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07581__S1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12786__17 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__inv_2
XFILLER_0_8_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09143_ net465 _03553_ _04061_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10655__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09074_ _03702_ _03722_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08025_ final_design.cpu.reg_window\[147\] final_design.cpu.reg_window\[179\] net825
+ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold720 final_design.cpu.reg_window\[938\] vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 final_design.cpu.reg_window\[798\] vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1228_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold742 final_design.cpu.reg_window\[761\] vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 final_design.cpu.reg_window\[872\] vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12534__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold764 final_design.cpu.reg_window\[232\] vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11742__A0 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout590_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 final_design.cpu.reg_window\[745\] vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__C1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 final_design.cpu.reg_window\[286\] vssd1 vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07410__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold797 final_design.cpu.reg_window\[351\] vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06844__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ _03358_ _04720_ _03565_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1016_X net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08927_ _03869_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout855_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09163__A1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08858_ net632 _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__nor2_1
XANTENNA__08910__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07809_ final_design.cpu.reg_window\[537\] final_design.cpu.reg_window\[569\] net863
+ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08789_ _03683_ _03686_ _03736_ _03739_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11425__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10820_ _01362_ _03909_ net1070 vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10751_ net74 _05466_ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_49_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout908_X net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13011__RESET_B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13470_ clknet_leaf_22_clk _00701_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[458\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10682_ _05421_ _05422_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ _06244_ net501 net340 net2020 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__a22o_1
XANTENNA__12222__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10565__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07324__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12352_ net2518 net363 net359 _06018_ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11981__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ net667 _03896_ net739 vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_75_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12283_ net570 _06213_ net506 net368 net1929 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_75_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14022_ clknet_leaf_171_clk _01253_ net1080 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1010\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12525__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ net739 _03965_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ net816 _05846_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__nor2_1
XANTENNA__07085__S net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input37_X net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ _05026_ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__inv_2
X_11096_ net2540 net1046 _05816_ _05817_ vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__a22o_1
XANTENNA__12289__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10047_ _04577_ _04598_ _04925_ _04965_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__a211oi_1
XANTENNA__13852__RESET_B net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 final_design.VGA_data_control.data_to_VGA\[18\] vssd1 vssd1 vccd1 vccd1 net1433
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_160_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold91 net146 vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11843__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13806_ clknet_leaf_120_clk _01037_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[794\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11998_ _06200_ net279 net400 net2313 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__a22o_1
XANTENNA__07114__A _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13737_ clknet_leaf_86_clk _00968_ net1235 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[725\]
+ sky130_fd_sc_hd__dfrtp_1
X_10949_ net84 net1060 vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07468__B2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11264__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10472__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13668_ clknet_leaf_94_clk _00899_ net1227 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[656\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12619_ net2475 final_design.reqhand.data_from_UART\[5\] _05080_ vssd1 vssd1 vccd1
+ vccd1 _01312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12213__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12166__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13599_ clknet_leaf_133_clk _00830_ net1166 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[587\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11972__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12516__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07784__A net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11724__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09830_ _04182_ _04745_ _04746_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout507 net508 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout518 net519 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_4
XFILLER_0_120_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09761_ _04143_ _04157_ _03590_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__o21ai_1
X_06973_ net765 _01917_ net756 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09145__A1 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08712_ final_design.CPU_instr_adr\[26\] _01630_ vssd1 vssd1 vccd1 vccd1 _03663_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_174_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09692_ _03071_ _03102_ _04496_ _03581_ _03165_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a311o_1
X_08643_ _02903_ net262 _03592_ _03040_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout269_A _06237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08574_ final_design.cpu.reg_window\[320\] final_design.cpu.reg_window\[352\] net862
+ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07525_ _01540_ _02475_ _01541_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11255__A2 _05953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12452__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1080_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_61_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout436_A _05847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07456_ net762 _02400_ net756 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06407_ final_design.CPU_instr_adr\[18\] vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07387_ final_design.cpu.reg_window\[66\] final_design.cpu.reg_window\[98\] net946
+ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout603_A _03627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09126_ _03631_ _03647_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__nor2_4
XFILLER_0_161_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11963__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11768__X _06227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09057_ _02441_ net629 _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__or3_1
XFILLER_0_142_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12507__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08008_ _02955_ _02956_ _02957_ _02958_ net696 net703 vssd1 vssd1 vccd1 vccd1 _02959_
+ sky130_fd_sc_hd__mux4_1
Xhold550 final_design.cpu.reg_window\[784\] vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 final_design.cpu.reg_window\[579\] vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold572 final_design.cpu.reg_window\[742\] vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09384__A1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold583 final_design.cpu.reg_window\[400\] vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11647__C net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 final_design.cpu.reg_window\[656\] vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11191__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ net450 _04877_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_142_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ clknet_leaf_48_clk _00208_ net1154 vssd1 vssd1 vccd1 vccd1 final_design.uart.bits_received\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09687__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07633__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__B net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11921_ net681 _06118_ _06124_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__or3_1
XFILLER_0_135_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07793__S1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11852_ _06102_ net282 net520 net2213 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10803_ net814 _05535_ _05537_ net974 vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__o22a_1
XANTENNA__11246__A2 _05943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12443__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11783_ net2325 net413 net287 _05935_ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_52_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13522_ clknet_leaf_26_clk _00753_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[510\]
+ sky130_fd_sc_hd__dfrtp_1
X_10734_ _01364_ _03940_ net1070 vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13453_ clknet_leaf_141_clk _00684_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[441\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10665_ _04677_ net254 _04990_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_149_Left_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12404_ _06102_ net347 net339 net2194 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__a22o_1
X_14245__1310 vssd1 vssd1 vccd1 vccd1 _14245__1310/HI net1310 sky130_fd_sc_hd__conb_1
XFILLER_0_134_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09072__B1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13384_ clknet_leaf_119_clk _00615_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[372\]
+ sky130_fd_sc_hd__dfrtp_1
X_10596_ final_design.CPU_instr_adr\[7\] _05239_ _05338_ _01371_ vssd1 vssd1 vccd1
+ vccd1 _05341_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10757__B2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11954__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07622__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12335_ net2521 net362 net353 _05891_ vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11001__A1_N net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12266_ _06196_ net515 net370 net2478 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__a22o_1
XANTENNA__06712__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11706__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14005_ clknet_leaf_26_clk _01236_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[993\]
+ sky130_fd_sc_hd__dfrtp_1
X_11217_ net669 _03976_ net745 vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a21o_1
XANTENNA__09308__B net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12197_ net231 net2361 net378 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__mux2_1
XANTENNA__11182__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07109__A final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11148_ _05855_ _05861_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_158_Left_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11079_ _05765_ _05779_ _05800_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__a21o_1
XANTENNA__12131__A0 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11065__S net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09395__A2_N _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12434__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12986__RESET_B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07310_ final_design.cpu.reg_window\[517\] final_design.cpu.reg_window\[549\] net904
+ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__mux2_1
XANTENNA__07536__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08290_ final_design.cpu.reg_window\[201\] final_design.cpu.reg_window\[233\] net842
+ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_167_Left_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07241_ _02188_ _02189_ _02190_ _02191_ net777 net791 vssd1 vssd1 vccd1 vccd1 _02192_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12198__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07172_ final_design.cpu.reg_window\[522\] final_design.cpu.reg_window\[554\] net919
+ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11945__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout304 net306 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__buf_4
Xfanout315 _05851_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_6
Xfanout326 _06285_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07019__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09813_ net543 net541 net540 net539 net453 net462 vssd1 vssd1 vccd1 vccd1 _04732_
+ sky130_fd_sc_hd__mux4_1
Xfanout337 net338 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__buf_6
XANTENNA__07916__A2 _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout348 net352 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_4
XANTENNA__10920__A1 _04550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout359 _06277_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__buf_4
XANTENNA_fanout386_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09744_ net545 net544 net543 net541 net453 net462 vssd1 vssd1 vccd1 vccd1 _04663_
+ sky130_fd_sc_hd__mux4_1
X_06956_ _01901_ _01906_ net758 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__mux2_1
XANTENNA__07453__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11483__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09675_ _04592_ _04593_ _04590_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12673__B2 final_design.data_from_mem\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_A _01784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06887_ final_design.cpu.reg_window\[851\] final_design.cpu.reg_window\[883\] net911
+ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08341__A2 _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ _03231_ _03576_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11770__Y _06228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11228__A2 _05930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ final_design.cpu.reg_window\[641\] final_design.cpu.reg_window\[673\] net854
+ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout720_A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_X net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk
+ sky130_fd_sc_hd__clkbuf_8
X_07508_ _01884_ _02457_ _01882_ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08284__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11930__C net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08488_ final_design.cpu.reg_window\[835\] final_design.cpu.reg_window\[867\] net863
+ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07439_ net897 _02382_ _02388_ _02375_ _02376_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__a32o_4
XTAP_TAPCELL_ROW_21_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10450_ _02763_ net602 vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_94_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11936__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09109_ net628 _04028_ _04029_ _02428_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10381_ net25 net1038 net1021 final_design.data_from_mem\[30\] vssd1 vssd1 vccd1
+ vccd1 _00134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12120_ net2224 net188 net390 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__mux2_1
XANTENNA__07628__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09409__A _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout975_X net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12051_ net2182 net190 net398 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold380 net156 vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09128__B _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 final_design.cpu.reg_window\[974\] vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12361__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11164__B2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ net677 _05714_ _05727_ net978 _05726_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__o221a_1
XANTENNA__13444__RESET_B net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10989__S net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09109__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 net877 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_2
Xfanout871 net876 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_2
Xfanout882 net883 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08459__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout893 _01687_ vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__buf_4
XFILLER_0_172_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07363__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ clknet_leaf_55_clk _00191_ net1160 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_4
Xhold1080 final_design.cpu.reg_window\[628\] vssd1 vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1091 final_design.cpu.reg_window\[123\] vssd1 vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07766__S1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11904_ _06003_ net2226 net274 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ clknet_leaf_87_clk _00122_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_29_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ net191 net1932 net268 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__mux2_1
XANTENNA__12416__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09150__Y _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08194__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11766_ net178 net2139 net417 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ clknet_leaf_162_clk _00736_ net1109 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[493\]
+ sky130_fd_sc_hd__dfrtp_1
X_10717_ net676 _05444_ _05455_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11697_ net209 net634 vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13436_ clknet_leaf_147_clk _00667_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[424\]
+ sky130_fd_sc_hd__dfrtp_1
X_10648_ net69 final_design.VGA_adr\[8\] vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__xor2_1
XANTENNA__09596__A1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12444__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13367_ clknet_leaf_141_clk _00598_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[355\]
+ sky130_fd_sc_hd__dfrtp_1
X_10579_ net64 _05324_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__and2_1
X_12318_ net1858 net196 net366 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__mux2_1
XANTENNA__09319__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11568__B net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13298_ clknet_leaf_27_clk _00529_ net1139 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[286\]
+ sky130_fd_sc_hd__dfrtp_1
X_12249_ net566 _06178_ net505 net372 net1520 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__a32o_1
XFILLER_0_139_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12352__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07454__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ final_design.cpu.reg_window\[149\] final_design.cpu.reg_window\[181\] net965
+ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__mux2_1
XANTENNA__08369__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07790_ final_design.cpu.reg_window\[281\] final_design.cpu.reg_window\[313\] net863
+ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__mux2_1
XANTENNA__06678__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08308__C1 _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06741_ net556 _01690_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12655__B2 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ net321 _04373_ _04378_ net319 _04375_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__a221o_1
X_06672_ final_design.cpu.reg_window\[666\] final_design.cpu.reg_window\[698\] net952
+ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08411_ final_design.cpu.reg_window\[261\] final_design.cpu.reg_window\[293\] net822
+ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__mux2_1
X_09391_ net483 _04309_ _04306_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11523__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_16_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08342_ _03290_ _03292_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__nor2_1
XANTENNA__09284__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__A1 _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09823__A2 _04153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08273_ net890 _03223_ _03212_ _03206_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__07834__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11630__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07224_ final_design.cpu.reg_window\[520\] final_design.cpu.reg_window\[552\] net920
+ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07155_ _02102_ _02103_ _02104_ _02105_ net782 net792 vssd1 vssd1 vccd1 vccd1 _02106_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout301_A net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__B2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07448__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11478__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ final_design.cpu.reg_window\[396\] final_design.cpu.reg_window\[428\] net927
+ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11146__A1 final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12343__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout768_A _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11494__A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07996__S1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 net179 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout189 _06045_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_2
X_07988_ final_design.cpu.reg_window\[272\] final_design.cpu.reg_window\[304\] net878
+ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__mux2_1
XANTENNA__07183__S net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ _04644_ _04645_ net480 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06939_ final_design.cpu.reg_window\[81\] final_design.cpu.reg_window\[113\] net911
+ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09658_ _04576_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07911__S net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08609_ _03559_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10397__X _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ _03134_ _04506_ _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__a21o_2
XANTENNA__11433__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11620_ net575 net421 _06167_ net299 net1498 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__a32o_1
XANTENNA__10409__B1 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ net574 net421 _06131_ net303 net1946 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10502_ net93 final_design.VGA_adr\[1\] vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_163_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire535 _02266_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_4
X_11482_ net193 net2457 net308 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire557 _01686_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13221_ clknet_leaf_4_clk _00452_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[209\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10433_ net1436 net1047 _05200_ net248 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_150_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13696__RESET_B net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12264__S net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__A1 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07358__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input64_A mem_adr_start[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ clknet_leaf_36_clk _00383_ net1134 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[140\]
+ sky130_fd_sc_hd__dfrtp_1
X_10364_ net6 net1037 net1020 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1 vccd1
+ _00117_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12103_ net2344 net219 net389 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ clknet_leaf_156_clk _00314_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_10295_ final_design.VGA_data_control.h_count\[2\] _05148_ vssd1 vssd1 vccd1 vccd1
+ _05149_ sky130_fd_sc_hd__and2b_1
XANTENNA__11137__A1 final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12334__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12034_ net2164 net244 net398 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__mux2_1
XANTENNA__07436__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11688__A2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout690 net698 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__buf_4
X_13985_ clknet_leaf_158_clk _01216_ net1113 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[973\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12637__B2 final_design.data_from_mem\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12936_ clknet_leaf_67_clk _00174_ net1223 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_8__f_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12867_ clknet_leaf_72_clk _00105_ net1245 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_122_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12439__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10748__A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11860__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11818_ net245 net2408 net266 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08164__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ net210 net2285 net417 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__mux2_1
XANTENNA__11612__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09281__A3 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06961__A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13419_ clknet_leaf_23_clk _00650_ net1157 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[407\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12174__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11376__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08241__B2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08960_ net630 _03898_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_5_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08888__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ _02856_ _02861_ net718 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__mux2_1
X_08891_ net259 _03837_ net1029 vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__a21oi_1
X_07842_ final_design.cpu.reg_window\[597\] final_design.cpu.reg_window\[629\] net884
+ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10351__A2 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07773_ _02720_ _02721_ _02722_ _02723_ net693 net712 vssd1 vssd1 vccd1 vccd1 _02724_
+ sky130_fd_sc_hd__mux4_1
X_09512_ _02965_ _03028_ _04351_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__and3_1
X_06724_ final_design.cpu.reg_window\[984\] final_design.cpu.reg_window\[1016\] net950
+ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14154__RESET_B net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ net465 _04079_ _04081_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__and3_1
X_06655_ _01602_ _01603_ _01604_ _01605_ net787 net804 vssd1 vssd1 vccd1 vccd1 _01606_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_82_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10658__A net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11851__A2 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout349_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09374_ net465 _04103_ _04257_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__and3_1
X_06586_ final_design.reqhand.instruction\[29\] final_design.data_from_mem\[29\] net985
+ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__mux2_4
XFILLER_0_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08325_ final_design.cpu.reg_window\[840\] final_design.cpu.reg_window\[872\] net861
+ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1160_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10811__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08256_ final_design.cpu.reg_window\[74\] final_design.cpu.reg_window\[106\] net852
+ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07207_ _02155_ _02157_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout304_X net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ final_design.cpu.reg_window\[462\] final_design.cpu.reg_window\[494\] net853
+ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11367__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1046_X net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_104_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07138_ _02085_ _02086_ _02087_ _02088_ net783 net793 vssd1 vssd1 vccd1 vccd1 _02089_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout885_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13036__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07069_ final_design.cpu.reg_window\[845\] final_design.cpu.reg_window\[877\] net916
+ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10080_ final_design.VGA_data_control.v_count\[2\] final_design.VGA_data_control.v_count\[1\]
+ final_design.VGA_data_control.v_count\[3\] vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07418__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06810__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11428__S net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08535__A2 _03481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09406__B _04324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09732__B2 _04341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07207__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12619__A1 final_design.reqhand.data_from_UART\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_113_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13770_ clknet_leaf_0_clk _01001_ net1078 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[758\]
+ sky130_fd_sc_hd__dfrtp_1
X_10982_ net53 _05708_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09496__B1 _04414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12721_ final_design.VGA_data_control.v_count\[2\] _06359_ vssd1 vssd1 vccd1 vccd1
+ _06362_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09422__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_154_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ _06313_ net1429 net992 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11055__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ net817 _02359_ _02392_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__or3b_1
XFILLER_0_33_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ net1489 net1012 net998 final_design.data_from_mem\[1\] vssd1 vssd1 vccd1
+ vccd1 _01276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_169_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11534_ net1532 net178 net525 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14253_ net1318 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11465_ net216 net2388 net308 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__mux2_1
XANTENNA__11358__A1 net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07088__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12555__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13204_ clknet_leaf_141_clk _00435_ net1185 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[192\]
+ sky130_fd_sc_hd__dfrtp_1
X_10416_ net1573 net1044 _05191_ net247 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__a22o_1
X_14184_ clknet_leaf_72_clk final_design.VGA_data_control.next_state\[0\] net1245
+ vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.state\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11396_ _04248_ net664 _06080_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__a21boi_4
XTAP_TAPCELL_ROW_78_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13135_ clknet_leaf_92_clk _00366_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[123\]
+ sky130_fd_sc_hd__dfrtp_1
X_10347_ wb_manage.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__and2_2
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13066_ clknet_leaf_1_clk _00297_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_10278_ final_design.uart.BAUD_counter\[27\] final_design.uart.BAUD_counter\[28\]
+ _05133_ final_design.uart.BAUD_counter\[29\] vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__a31o_1
XANTENNA__08501__A _02330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09184__C1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12017_ _06219_ net288 net402 net2190 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__a22o_1
XANTENNA__09723__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11530__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13968_ clknet_leaf_111_clk _01199_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[956\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11294__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12169__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12919_ clknet_leaf_90_clk _00157_ net1232 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dfrtp_1
X_13899_ clknet_leaf_19_clk _01130_ net1122 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[887\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06440_ wb_manage.BUSY_O net34 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11597__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08110_ final_design.cpu.reg_window\[588\] final_design.cpu.reg_window\[620\] net847
+ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09090_ _03708_ _03720_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08041_ _01853_ net617 vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11349__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12546__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold902 final_design.cpu.reg_window\[510\] vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 final_design.cpu.reg_window\[331\] vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12010__A2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold924 final_design.cpu.reg_window\[580\] vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 final_design.cpu.reg_window\[127\] vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold946 final_design.cpu.reg_window\[104\] vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 net169 vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 final_design.cpu.reg_window\[757\] vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ net264 _04908_ _04910_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__and3_1
Xhold979 final_design.cpu.reg_window\[355\] vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
X_08943_ _02462_ _03883_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout299_A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ final_design.CPU_instr_adr\[29\] net1030 _03819_ _03822_ vssd1 vssd1 vccd1
+ vccd1 _00240_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07825_ final_design.cpu.reg_window\[85\] final_design.cpu.reg_window\[117\] net884
+ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11772__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07756_ _01690_ net621 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__or2_1
XANTENNA__08557__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06707_ net898 _01650_ _01656_ _01643_ _01644_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__a32o_2
XFILLER_0_17_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07687_ _02637_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout254_X net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_A _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09426_ _02899_ net443 net439 _02898_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06638_ net765 _01588_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09357_ net490 _04275_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13970__RESET_B net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06569_ _01516_ _01517_ _01518_ _01519_ net788 net806 vssd1 vssd1 vccd1 vccd1 _01520_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1163_X net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08989__C1 _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08308_ net605 _03257_ _03232_ _02155_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__o211a_1
XFILLER_0_164_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08145__X _03096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09288_ net614 _03550_ _03524_ net561 vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08239_ _03186_ _03187_ _03188_ _03189_ net691 net702 vssd1 vssd1 vccd1 vccd1 _03190_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12537__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11012__A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11250_ net428 net580 _05952_ net316 net1604 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__a32o_1
XFILLER_0_127_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12001__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout888_X net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ _05088_ _05089_ _00039_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_56_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13000__Q final_design.CPU_instr_adr\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ net432 net584 _05891_ net317 net2398 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__a32o_1
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06767__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07636__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ net2573 _04997_ _05036_ _01404_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_state\[1\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06862__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10063_ _04290_ _04328_ _04389_ _04981_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__and4_1
XANTENNA__09136__B _04053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08064__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11512__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07716__B1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14005__RESET_B net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13822_ clknet_leaf_147_clk _01053_ net1127 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[810\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10079__A1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07371__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13753_ clknet_leaf_168_clk _00984_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[741\]
+ sky130_fd_sc_hd__dfrtp_1
X_10965_ _05692_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12704_ _06340_ _06344_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__or2_1
X_13684_ clknet_leaf_104_clk _00915_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[672\]
+ sky130_fd_sc_hd__dfrtp_1
X_10896_ net2523 net1043 _05624_ _05626_ vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12635_ final_design.VGA_data_control.ready_data\[5\] net1035 net990 final_design.data_from_mem\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_130_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11579__A1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12566_ final_design.uart.receiving final_design.uart.working_data\[3\] vssd1 vssd1
+ vccd1 vccd1 _06288_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06715__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11517_ net2341 net205 net524 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ net597 _06158_ _06260_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_117_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12528__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14236_ net1301 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
Xhold209 final_design.cpu.reg_window\[685\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ net242 net647 vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_169_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08747__A2 _01598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14167_ clknet_leaf_78_clk _01341_ net1250 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12452__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ _04420_ net664 vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__nand2_1
XANTENNA__07546__S net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ clknet_leaf_21_clk _00349_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11576__B net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14098_ clknet_leaf_71_clk _01295_ net1243 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_13049_ clknet_leaf_166_clk _00280_ net1082 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11503__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07610_ final_design.cpu.reg_window\[733\] final_design.cpu.reg_window\[765\] net880
+ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__mux2_1
XANTENNA__11592__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08590_ _03537_ _03538_ _03539_ _03540_ net694 net713 vssd1 vssd1 vccd1 vccd1 _03541_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_3_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06930__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06930__B2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07541_ final_design.cpu.reg_window\[991\] final_design.cpu.reg_window\[1023\] net923
+ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
XANTENNA__11806__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09475__A3 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07472_ _02420_ _02421_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__or2_2
XFILLER_0_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09211_ _02800_ _02834_ _02802_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_174_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06423_ final_design.reqhand.instruction\[5\] vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
XANTENNA__10490__B2 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11531__S net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09142_ net614 _03549_ net531 _02422_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12231__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09073_ _02242_ _02436_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13310__RESET_B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout214_A _05941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08024_ final_design.cpu.reg_window\[211\] final_design.cpu.reg_window\[243\] net825
+ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold710 final_design.cpu.reg_window\[159\] vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold721 final_design.cpu.reg_window\[587\] vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 final_design.cpu.reg_window\[952\] vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold743 final_design.cpu.reg_window\[583\] vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold754 final_design.cpu.reg_window\[706\] vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 final_design.cpu.reg_window\[870\] vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1123_A net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 final_design.cpu.reg_window\[881\] vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 final_design.cpu.reg_window\[841\] vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11486__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07410__A2 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09975_ _04221_ _04533_ _04539_ _04728_ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a221o_1
Xhold798 final_design.cpu.reg_window\[144\] vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06844__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout583_A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ _03797_ _03868_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_51_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09699__A0 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ _03658_ _03778_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout750_A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout848_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08795__B _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07808_ final_design.cpu.reg_window\[601\] final_design.cpu.reg_window\[633\] net859
+ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__mux2_1
X_08788_ _03679_ _03680_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__nor2_1
XANTENNA__06596__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11258__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07739_ final_design.cpu.reg_window\[922\] final_design.cpu.reg_window\[954\] net872
+ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _05485_ _05486_ _05466_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_49_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09409_ _04325_ _04326_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10681_ _05402_ _05404_ _05400_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07882__C1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11441__S net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12420_ _06024_ net563 net500 net339 net1920 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__a32o_1
XFILLER_0_164_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_7__f_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_97_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12351_ _06235_ net503 net362 final_design.cpu.reg_window\[820\] vssd1 vssd1 vccd1
+ vccd1 _01063_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06988__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11302_ final_design.data_from_mem\[19\] net235 net233 vssd1 vssd1 vccd1 vccd1 _05998_
+ sky130_fd_sc_hd__a21o_2
XANTENNA__06988__B2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12282_ net566 _06212_ net505 net368 net1780 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_75_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14021_ clknet_leaf_150_clk _01252_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1009\]
+ sky130_fd_sc_hd__dfrtp_1
X_11233_ net669 _03962_ net743 vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11164_ net2466 net317 _05876_ net434 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ final_design.VGA_data_control.v_count\[5\] net1064 _05023_ vssd1 vssd1 vccd1
+ vccd1 _05026_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_164_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11095_ _05798_ _05815_ net1016 vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__o21a_1
X_10046_ net736 _04576_ _04597_ _04421_ _04423_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a32o_1
XFILLER_0_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_160_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 final_design.VGA_data_control.data_to_VGA\[19\] vssd1 vssd1 vccd1 vccd1 net1423
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 final_design.cpu.reg_window\[716\] vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 net155 vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09153__Y _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13805_ clknet_leaf_127_clk _01036_ net1193 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[793\]
+ sky130_fd_sc_hd__dfrtp_1
X_11997_ _06199_ net278 net400 net2251 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07114__B _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ _05634_ _05653_ _05675_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__a21o_1
X_13736_ clknet_leaf_118_clk _00967_ net1195 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[724\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10472__A1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09610__A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10879_ net81 net1055 vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__nor2_2
XANTENNA__10756__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ clknet_leaf_1_clk _00898_ net1077 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[655\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12447__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12618_ final_design.uart.working_data\[5\] net1512 _05080_ vssd1 vssd1 vccd1 vccd1
+ _01311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13598_ clknet_leaf_18_clk _00829_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[586\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12549_ _06212_ net343 net323 net2033 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14219_ net1288 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XANTENNA__12182__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11724__A1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout508 net513 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__buf_2
Xfanout519 _06259_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_4
X_09760_ _04659_ _04677_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__nand2_1
X_06972_ net773 _01922_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__or2_2
XANTENNA__08628__A_N net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08711_ final_design.CPU_instr_adr\[26\] _01630_ vssd1 vssd1 vccd1 vccd1 _03662_
+ sky130_fd_sc_hd__nand2_1
X_09691_ _04340_ _04608_ _04609_ _04604_ _04605_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a311o_1
XFILLER_0_174_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11526__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1090 net1095 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__buf_2
X_08642_ _02838_ _02901_ _03030_ _03591_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__and4_1
X_08573_ _02424_ net613 vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__nand2_2
X_07524_ _01567_ _01570_ _02474_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08656__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09853__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07455_ net772 _02405_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10463__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11660__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout331_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1073_A final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout429_A net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06406_ final_design.CPU_instr_adr\[24\] vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07386_ _02333_ _02334_ _02335_ _02336_ net785 net803 vssd1 vssd1 vccd1 vccd1 _02337_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12204__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09125_ net971 net969 net975 vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09056_ _02439_ _02440_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout798_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ final_design.cpu.reg_window\[528\] final_design.cpu.reg_window\[560\] net879
+ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold540 final_design.cpu.reg_window\[243\] vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold551 final_design.cpu.reg_window\[91\] vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_3_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07186__S net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 final_design.cpu.reg_window\[585\] vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 final_design.cpu.reg_window\[376\] vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold584 final_design.cpu.reg_window\[911\] vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold595 final_design.cpu.reg_window\[449\] vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout965_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_X net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_15__f_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_70_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09958_ _03488_ _04145_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ net90 net93 vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__xor2_1
XANTENNA__11436__S net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09687__A3 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11920_ net177 net2155 net274 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11851_ _06101_ net281 net520 net2308 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ net972 _05534_ _05536_ net968 vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ net2397 net413 net284 _05929_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10733_ _05469_ _05470_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__or2_1
X_13521_ clknet_leaf_108_clk _00752_ net1213 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[509\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ clknet_leaf_121_clk _00683_ net1198 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[440\]
+ sky130_fd_sc_hd__dfrtp_1
X_10664_ net1483 net1042 net1015 _05405_ vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__a22o_1
XANTENNA_input94_A memory_size[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12403_ _06101_ net347 net339 net2118 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13383_ clknet_leaf_16_clk _00614_ net1097 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[371\]
+ sky130_fd_sc_hd__dfrtp_1
X_10595_ net971 _05338_ _05339_ net969 vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__o22a_1
XFILLER_0_24_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11954__A1 _06155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12334_ _06230_ net502 net362 net2039 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07622__A2 _02570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12265_ net581 _06195_ net512 net369 net2231 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11706__A1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14004_ clknet_leaf_101_clk _01235_ net1188 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[992\]
+ sky130_fd_sc_hd__dfrtp_1
X_11216_ net2443 net315 _05922_ net427 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__a22o_1
X_12196_ net679 _06124_ _06262_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__or3_4
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11147_ final_design.reqhand.data_from_UART\[1\] final_design.data_from_mem\[1\]
+ net249 vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__mux2_1
XANTENNA__12730__S final_design.VGA_data_control.v_count\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10390__B1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07824__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11078_ _05763_ _05779_ _05782_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__a21bo_1
X_10029_ net497 _04836_ _04838_ _04231_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__a31o_1
XANTENNA__09989__B1_N _04409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11642__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13719_ clknet_leaf_143_clk _00950_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[707\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10445__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10486__A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12177__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07240_ final_design.cpu.reg_window\[7\] final_design.cpu.reg_window\[39\] net915
+ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12198__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07171_ final_design.cpu.reg_window\[586\] final_design.cpu.reg_window\[618\] net919
+ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__mux2_1
XANTENNA__08497__S0 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12955__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14179__RESET_B net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout305 net306 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11173__A2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout316 _05851_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_4
XANTENNA__12370__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_8
X_09812_ net492 _04368_ _04727_ _04730_ net263 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__o311a_1
Xfanout338 _06282_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_4
Xfanout349 net350 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10920__A2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06955_ _01902_ _01903_ _01904_ _01905_ net775 net791 vssd1 vssd1 vccd1 vccd1 _01906_
+ sky130_fd_sc_hd__mux4_1
X_09743_ net319 _04278_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout281_A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12122__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A _06271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ _02838_ _04352_ net322 _03035_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06886_ net767 _01836_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__nor2_1
X_08625_ _03262_ _03574_ _03573_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__o21bai_1
XANTENNA__11881__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1190_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A _01966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08556_ final_design.cpu.reg_window\[705\] final_design.cpu.reg_window\[737\] net851
+ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12425__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__C _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06874__A _01815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07507_ _01884_ _02457_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08487_ net722 _03431_ net731 vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout713_A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07438_ net897 _02382_ _02388_ _02375_ _02376_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__a32oi_1
XTAP_TAPCELL_ROW_21_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12189__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout501_X net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07369_ final_design.cpu.reg_window\[643\] final_design.cpu.reg_window\[675\] net942
+ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09054__B2 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ _02426_ _02427_ net628 vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__a21oi_1
X_10380_ net23 net1036 net1019 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1
+ vccd1 _00133_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_131_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ _02159_ _02443_ _02130_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12050_ net2323 net192 net396 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__mux2_1
Xhold370 final_design.cpu.reg_window\[660\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 final_design.reqhand.instruction\[14\] vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ net1067 _05724_ _05239_ final_design.CPU_instr_adr\[26\] vssd1 vssd1 vccd1
+ vccd1 _05727_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout968_X net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold392 final_design.cpu.reg_window\[203\] vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11164__A2 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout850 net851 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
Xfanout861 net864 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_4
Xfanout872 net875 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__clkbuf_4
Xfanout883 net886 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_4
Xfanout894 _01437_ vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_172_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12952_ clknet_leaf_55_clk _00190_ net1160 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_4
Xhold1070 final_design.cpu.reg_window\[882\] vssd1 vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 final_design.cpu.reg_window\[353\] vssd1 vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10675__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ net202 net1975 net274 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__mux2_1
Xhold1092 final_design.cpu.reg_window\[319\] vssd1 vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10675__B2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13413__RESET_B net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ clknet_leaf_88_clk _00121_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11834_ net193 net2407 net267 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__mux2_1
XANTENNA__12416__A2 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11765_ net181 net2123 net419 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__mux2_1
XANTENNA__11624__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ net814 _05452_ _05454_ net974 vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__o22a_1
X_13504_ clknet_leaf_35_clk _00735_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[492\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input97_X net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11696_ net428 net579 _06206_ net296 net1711 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__a32o_1
XFILLER_0_165_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ _05354_ _05374_ _05373_ _05371_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13435_ clknet_leaf_153_clk _00666_ net1117 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[423\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11927__B2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13366_ clknet_leaf_126_clk _00597_ net1192 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[354\]
+ sky130_fd_sc_hd__dfrtp_1
X_10578_ net677 _05310_ _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__o21a_1
XANTENNA__08504__A _02325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12317_ net1770 net198 net366 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__mux2_1
XANTENNA__09319__B net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13297_ clknet_leaf_111_clk _00528_ net1214 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[285\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09348__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12248_ net571 _06177_ net506 net372 net1580 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__a32o_1
XFILLER_0_139_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11865__A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ net1696 net205 net380 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__mux2_1
XANTENNA__12460__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07454__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__B net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_13 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06678__B _01628_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ _01499_ net672 _01689_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__or3b_1
XFILLER_0_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08859__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06671_ final_design.cpu.reg_window\[730\] final_design.cpu.reg_window\[762\] net953
+ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08410_ final_design.cpu.reg_window\[325\] final_design.cpu.reg_window\[357\] net822
+ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__mux2_1
X_09390_ _04307_ _04308_ net478 vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__mux2_2
XANTENNA__08385__S net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12407__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08341_ net605 _03287_ _03263_ _02184_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10418__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10969__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08272_ _03217_ _03222_ net718 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07223_ final_design.cpu.reg_window\[584\] final_design.cpu.reg_window\[616\] net920
+ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07729__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07154_ final_design.cpu.reg_window\[266\] final_design.cpu.reg_window\[298\] net936
+ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__mux2_1
XANTENNA__08244__C1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06633__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__A2 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12591__B2 final_design.data_from_mem\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07085_ final_design.cpu.reg_window\[460\] final_design.cpu.reg_window\[492\] net929
+ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1036_A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13995__RESET_B net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11146__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout496_A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__S net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__B1 _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1203_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11494__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07987_ final_design.cpu.reg_window\[336\] final_design.cpu.reg_window\[368\] net878
+ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__mux2_1
Xfanout179 _06081_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_2
XANTENNA_fanout663_A _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06938_ _01885_ _01886_ _01887_ _01888_ net778 net791 vssd1 vssd1 vccd1 vccd1 _01889_
+ sky130_fd_sc_hd__mux4_1
X_09726_ net560 net559 net558 net556 net455 net464 vssd1 vssd1 vccd1 vccd1 _04645_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_87_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10657__A1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ _04190_ _04575_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__and2_1
XANTENNA__10657__B2 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06869_ _01464_ _01468_ _01475_ _01483_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__or4_4
XANTENNA_fanout830_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11854__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout928_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _02356_ net481 vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__or2_1
XANTENNA__08295__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09588_ _03134_ _04506_ net451 vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10409__B2 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08539_ final_design.cpu.reg_window\[257\] final_design.cpu.reg_window\[289\] net849
+ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ net237 net642 vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_61_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ net734 _04825_ net252 _04990_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_107_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11481_ net194 net2324 net307 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11302__X _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire558 _01657_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_4
X_13220_ clknet_leaf_106_clk _00451_ net1227 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[208\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07639__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ net601 _02961_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_150_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07133__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07589__A1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12582__B2 final_design.data_from_mem\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ clknet_leaf_134_clk _00382_ net1165 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[139\]
+ sky130_fd_sc_hd__dfrtp_1
X_10363_ net5 net1036 net1019 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1
+ _00116_ sky130_fd_sc_hd__o22a_1
X_12102_ net2096 net244 net390 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09707__X _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13082_ clknet_leaf_164_clk _00313_ net1108 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input57_A mem_adr_start[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ final_design.VGA_data_control.data_to_VGA\[7\] final_design.VGA_data_control.data_to_VGA\[6\]
+ final_design.VGA_data_control.h_count\[1\] vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__mux2_1
XANTENNA__11137__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12033_ net2009 net237 net396 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__mux2_1
XANTENNA__07436__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09750__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout680 _02329_ vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_2
Xfanout691 net698 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_8
X_13984_ clknet_leaf_38_clk _01215_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[972\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ clknet_leaf_68_clk _00173_ net1221 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12866_ clknet_leaf_72_clk _00104_ net1245 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_122_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ net238 net2216 net267 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12270__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07816__A2 _02763_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11748_ net212 net2204 net416 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07372__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12455__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ net240 net636 vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13418_ clknet_leaf_2_clk _00649_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[406\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12022__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13349_ clknet_leaf_150_clk _00580_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[337\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12190__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ _02857_ _02858_ _02859_ _02860_ net684 net699 vssd1 vssd1 vccd1 vccd1 _02861_
+ sky130_fd_sc_hd__mux4_1
X_08890_ final_design.CPU_instr_adr\[27\] _03799_ vssd1 vssd1 vccd1 vccd1 _03837_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10336__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ final_design.cpu.reg_window\[661\] final_design.cpu.reg_window\[693\] net886
+ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__mux2_1
X_07772_ final_design.cpu.reg_window\[920\] final_design.cpu.reg_window\[952\] net869
+ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__mux2_1
XANTENNA__12089__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10004__A _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10639__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06723_ net762 _01673_ net756 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__o21a_1
XANTENNA__11836__A0 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09511_ _02965_ _04351_ _03028_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11534__S net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06938__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ _02769_ _03597_ _04046_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__o21a_1
X_06654_ final_design.cpu.reg_window\[410\] final_design.cpu.reg_window\[442\] net953
+ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__mux2_1
XANTENNA__06628__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _03606_ _04046_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__nand2_1
X_06585_ net900 _01528_ _01534_ _01521_ _01522_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__a32o_2
XANTENNA__12970__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_A _05910_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11064__A1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08324_ net718 _03268_ net730 vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__o21a_1
XANTENNA__12261__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10945__Y _05673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08255_ net720 _03205_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10811__B2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12365__S net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1153_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07206_ net673 _01537_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12013__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08186_ final_design.cpu.reg_window\[270\] final_design.cpu.reg_window\[302\] net852
+ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07137_ final_design.cpu.reg_window\[523\] final_design.cpu.reg_window\[555\] net937
+ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1039_X net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07440__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ _02015_ _02016_ _02017_ _02018_ net777 net797 vssd1 vssd1 vccd1 vccd1 _02019_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout780_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12316__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10327__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07418__S1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07194__S net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13076__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13005__RESET_B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07207__B _02157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07922__S net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ _03068_ _04627_ _03101_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a21oi_1
X_10981_ net813 _05704_ _05707_ _05696_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12720_ _06355_ _06356_ _06360_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12651_ final_design.VGA_data_control.ready_data\[13\] net1032 net988 final_design.data_from_mem\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__a22o_1
XANTENNA__09248__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_0__f_clk_X clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11055__A1 _04325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11602_ net817 _02358_ net815 vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__and3b_4
XFILLER_0_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12582_ net1619 net1012 net998 final_design.data_from_mem\[0\] vssd1 vssd1 vccd1
+ vccd1 _01275_ sky130_fd_sc_hd__a22o_1
XANTENNA__12252__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07354__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10802__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10802__B2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11533_ net1722 net180 net527 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08471__A2 _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07369__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14252_ net1317 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_163_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11464_ net215 net646 vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__and2_1
XANTENNA__12004__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10415_ _03287_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13203_ clknet_leaf_34_clk _00434_ net1130 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[191\]
+ sky130_fd_sc_hd__dfrtp_1
X_14183_ clknet_leaf_56_clk _01357_ net1162 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11395_ net664 _06077_ _06079_ net599 vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__o31a_1
XANTENNA__13846__RESET_B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09437__X _04356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10346_ net1522 net1023 net1000 final_design.data_from_mem\[31\] vssd1 vssd1 vccd1
+ vccd1 _00103_ sky130_fd_sc_hd__a22o_1
X_13134_ clknet_leaf_115_clk _00365_ net1203 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12307__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ clknet_leaf_95_clk _00296_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[53\]
+ sky130_fd_sc_hd__dfrtp_1
X_10277_ net1541 _05134_ _05136_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__a21oi_1
X_12016_ _06218_ net290 net402 net2040 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09184__B1 _01536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13967_ clknet_leaf_89_clk _01198_ net1234 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[955\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12086__A3 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11294__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12918_ clknet_leaf_10_clk _00156_ net1091 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12491__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13898_ clknet_leaf_4_clk _01129_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[886\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12849_ clknet_leaf_78_clk _00087_ net1250 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11046__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11046__B2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12243__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06972__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11597__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08040_ net888 _02972_ _02978_ _02984_ _02990_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__o32a_4
XFILLER_0_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11349__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold903 final_design.cpu.reg_window\[357\] vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09411__A1 _04158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold914 final_design.cpu.reg_window\[758\] vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 final_design.cpu.reg_window\[636\] vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold936 final_design.cpu.reg_window\[484\] vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 final_design.cpu.reg_window\[101\] vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 final_design.cpu.reg_window\[818\] vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 final_design.cpu.reg_window\[258\] vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ _02738_ net447 net439 _02735_ _04909_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11529__S net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_11__f_clk_X clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ _01789_ _01790_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__nand2b_1
X_08873_ net260 _03821_ net1030 vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_32_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout194_A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07824_ final_design.cpu.reg_window\[149\] final_design.cpu.reg_window\[181\] net886
+ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__mux2_1
XANTENNA__07742__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11772__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11809__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07755_ _02670_ _02671_ _02701_ _02703_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__o22a_1
XANTENNA__12077__A3 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_A net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11285__A1 final_design.data_from_mem\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06706_ net899 _01650_ _01656_ _01643_ _01644_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__a32oi_2
X_07686_ net626 _02635_ _02636_ net562 vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__a211oi_2
XANTENNA__12482__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10021__X _04940_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07043__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09425_ _04342_ _04343_ _04339_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_94_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06637_ _01584_ _01585_ _01586_ _01587_ net789 net807 vssd1 vssd1 vccd1 vccd1 _01588_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout247_X net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout626_A _02513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12234__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ _04058_ _04060_ net478 vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__mux2_1
X_06568_ final_design.cpu.reg_window\[157\] final_design.cpu.reg_window\[189\] net959
+ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__mux2_1
XANTENNA__08438__C1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07336__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08307_ _02157_ net605 vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__and2_1
XANTENNA__12095__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09287_ _03418_ _04097_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__or3_1
XFILLER_0_173_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06499_ _01446_ _01447_ _01448_ _01449_ net779 net792 vssd1 vssd1 vccd1 vccd1 _01450_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1156_X net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800__31 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__inv_2
X_08238_ final_design.cpu.reg_window\[523\] final_design.cpu.reg_window\[555\] net856
+ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout995_A _06296_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08169_ final_design.cpu.reg_window\[975\] final_design.cpu.reg_window\[1007\] net826
+ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__mux2_1
X_10200_ net1065 net35 vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11180_ net656 net239 vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_56_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06821__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ final_design.VGA_data_control.v_count\[0\] _01399_ _05000_ _01401_ vssd1
+ vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_128_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11439__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08684__A_N _03617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _04249_ _04252_ _04356_ _04358_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__o22a_1
XANTENNA__09705__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08064__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07716__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09704__Y _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ clknet_leaf_13_clk _01052_ net1101 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[809\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12068__A3 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13752_ clknet_leaf_131_clk _00983_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[740\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12473__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10964_ _05689_ _05691_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07575__S0 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__X _04639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12703_ _06341_ _06343_ _06338_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__a21oi_2
XANTENNA__14045__RESET_B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13683_ clknet_leaf_36_clk _00914_ net1133 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[671\]
+ sky130_fd_sc_hd__dfrtp_1
X_10895_ _05606_ _05623_ _05625_ net1018 vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11902__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07888__A _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12634_ _06304_ net1547 net994 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__mux2_1
XANTENNA__12225__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09316__S1 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06792__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08483__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11579__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12565_ net1398 _06287_ _06286_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12240__A3 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11203__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11516_ net1996 net207 net525 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ _06156_ net349 net332 net2087 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14235_ net1300 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_150_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11447_ net229 net2503 net308 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__mux2_1
XANTENNA__10539__B1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14166_ clknet_leaf_78_clk _01340_ net1251 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_11378_ _01570_ net650 _06064_ _05853_ net664 vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a221o_1
XANTENNA__08071__X _03022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06731__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10329_ net1594 net1025 net1002 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1
+ vccd1 _00086_ sky130_fd_sc_hd__a22o_1
X_13117_ clknet_leaf_10_clk _00348_ net1092 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14097_ clknet_leaf_96_clk _01294_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09157__A0 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13048_ clknet_leaf_133_clk _00279_ net1166 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1250 net1251 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_1_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11592__B net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06930__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11267__A1 final_design.data_from_mem\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ final_design.cpu.reg_window\[799\] final_design.cpu.reg_window\[831\] net929
+ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07471_ _02420_ _02421_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11812__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06422_ final_design.data_from_mem\[4\] vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09210_ _02867_ _02897_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__nor2_1
XANTENNA__12216__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08393__S net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09141_ net537 net536 net534 net533 net461 _03518_ vssd1 vssd1 vccd1 vccd1 _04060_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08435__A2 _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09072_ _02242_ _02436_ net628 vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08023_ final_design.cpu.reg_window\[19\] final_design.cpu.reg_window\[51\] net825
+ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold700 final_design.cpu.reg_window\[772\] vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout207_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold711 final_design.cpu.reg_window\[417\] vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold722 final_design.cpu.reg_window\[161\] vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07737__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold733 final_design.cpu.reg_window\[456\] vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 final_design.cpu.reg_window\[473\] vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06641__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold755 final_design.cpu.reg_window\[175\] vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_153_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold766 final_design.cpu.reg_window\[916\] vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold777 final_design.cpu.reg_window\[38\] vssd1 vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 final_design.cpu.reg_window\[921\] vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 final_design.cpu.reg_window\[934\] vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ net490 _04487_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ final_design.CPU_instr_adr\[23\] _03796_ vssd1 vssd1 vccd1 vccd1 _03868_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_51_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09699__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_A _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__B net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ _01510_ _02476_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_168_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ final_design.cpu.reg_window\[665\] final_design.cpu.reg_window\[697\] net859
+ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__mux2_1
X_08787_ _03684_ _03737_ _03681_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout743_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11258__A1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__A_N _01750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ final_design.cpu.reg_window\[986\] final_design.cpu.reg_window\[1018\] net873
+ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout910_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07669_ final_design.cpu.reg_window\[158\] final_design.cpu.reg_window\[190\] net847
+ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_9_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09408_ _04325_ _04326_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__or2_1
X_10680_ _05418_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__nand2_1
XANTENNA__12207__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06816__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12758__B2 final_design.VGA_adr\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09339_ _04103_ _04257_ net465 vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12222__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12350_ _06234_ net500 net360 net2293 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__a22o_1
XANTENNA__13438__RESET_B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06988__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11301_ net425 net566 _05997_ net315 net1758 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__a32o_1
XANTENNA__11981__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12281_ net571 _06211_ net506 net368 net1749 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11232_ final_design.data_from_mem\[11\] _05914_ _05917_ vssd1 vssd1 vccd1 vccd1
+ _05936_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_75_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14020_ clknet_leaf_106_clk _01251_ net1206 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[1008\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11677__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ net657 net588 net241 vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_112_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09139__A0 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ net1064 _05023_ _05025_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_164_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11094_ _05798_ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_164_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12289__A3 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11693__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ _04632_ _04634_ _04421_ _04423_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10801__S net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08478__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 net167 vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07382__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold71 net111 vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07235__X _02186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold82 final_design.VGA_data_control.data_to_VGA\[25\] vssd1 vssd1 vccd1 vccd1 net1435
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 final_design.VGA_data_control.ready_data\[22\] vssd1 vssd1 vccd1 vccd1 net1446
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ clknet_leaf_121_clk _01035_ net1197 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[792\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11996_ _06198_ net288 net402 net2289 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__a22o_1
XANTENNA__08114__B2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13735_ clknet_leaf_9_clk _00966_ net1090 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[723\]
+ sky130_fd_sc_hd__dfrtp_1
X_10947_ _05632_ _05653_ _05652_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_156_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06676__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10472__A2 _04805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06726__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13666_ clknet_leaf_28_clk _00897_ net1141 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[654\]
+ sky130_fd_sc_hd__dfrtp_1
X_10878_ net81 net1056 vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_119_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07411__A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12617_ net2127 final_design.reqhand.data_from_UART\[3\] _05080_ vssd1 vssd1 vccd1
+ vccd1 _01310_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13861__RESET_B net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13597_ clknet_leaf_33_clk _00828_ net1129 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[585\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12213__A3 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12548_ _06211_ net346 net323 net2065 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11972__A2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13108__RESET_B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12463__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _06139_ net351 net332 net2054 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__a22o_1
XANTENNA_2 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12791__22 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__inv_2
XFILLER_0_50_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14218_ net1287 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08242__A _02097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14149_ clknet_leaf_80_clk _01323_ net1249 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09057__B net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout509 net513 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_4
X_06971_ _01918_ _01919_ _01920_ _01921_ net788 net806 vssd1 vssd1 vccd1 vccd1 _01922_
+ sky130_fd_sc_hd__mux4_1
X_08710_ _01359_ _01599_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__nand2_1
XANTENNA__08889__C1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ net492 _04338_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__nand2_1
Xfanout1080 net1104 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__buf_2
Xfanout1091 net1094 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_4
X_08641_ _03030_ _03591_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08572_ _02425_ net626 vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__nor2_2
XANTENNA__10012__A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07523_ _01601_ _02473_ _01571_ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__a21o_1
XFILLER_0_159_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07454_ _02401_ _02402_ _02403_ _02404_ net783 net802 vssd1 vssd1 vccd1 vccd1 _02405_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10463__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11660__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06405_ final_design.CPU_instr_adr\[26\] vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
XANTENNA__12935__Q net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07385_ final_design.cpu.reg_window\[386\] final_design.cpu.reg_window\[418\] net940
+ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout324_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1066_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ net1006 net1004 vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__nand2_1
XANTENNA__11412__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09947__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ _03725_ _03727_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11963__A2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12373__S net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1233_A net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07467__S net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08006_ final_design.cpu.reg_window\[592\] final_design.cpu.reg_window\[624\] net879
+ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold530 final_design.cpu.reg_window\[466\] vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout693_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold541 final_design.cpu.reg_window\[890\] vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold552 final_design.cpu.reg_window\[177\] vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold563 final_design.cpu.reg_window\[867\] vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 final_design.cpu.reg_window\[404\] vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A3 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold585 final_design.cpu.reg_window\[965\] vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 final_design.cpu.reg_window\[84\] vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09957_ _03557_ _04875_ _04874_ _03652_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout860_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _03798_ _03852_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__or2_1
X_09888_ net79 net734 _04805_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__or3_1
XANTENNA__07778__S0 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ final_design.CPU_instr_adr\[13\] final_design.CPU_instr_adr\[12\] _03789_
+ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11850_ _06100_ net279 net520 net2256 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__a22o_1
XANTENNA__12428__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10801_ final_design.CPU_instr_adr\[17\] _03919_ net1070 vssd1 vssd1 vccd1 vccd1
+ _05536_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ net2530 net412 _06231_ net433 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13520_ clknet_leaf_114_clk _00751_ net1211 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[508\]
+ sky130_fd_sc_hd__dfrtp_1
X_10732_ _05464_ _05468_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13451_ clknet_leaf_15_clk _00682_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[439\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10663_ _05402_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__xor2_1
X_12402_ _06100_ net344 net339 net1989 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__a22o_1
XANTENNA__07607__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input87_A memory_size[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10594_ final_design.CPU_instr_adr\[7\] _03995_ net1071 vssd1 vssd1 vccd1 vccd1 _05339_
+ sky130_fd_sc_hd__mux2_1
X_13382_ clknet_leaf_165_clk _00613_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[370\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11954__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12333_ _06229_ net503 net362 net2171 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12264_ net231 net2470 net370 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__mux2_1
XANTENNA__11706__A2 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14003_ clknet_leaf_35_clk _01234_ net1132 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[991\]
+ sky130_fd_sc_hd__dfrtp_1
X_11215_ net654 net575 net219 vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__and3_1
X_12195_ net1568 net176 net381 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__mux2_1
XANTENNA_input42_X net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11146_ final_design.CPU_instr_adr\[1\] net741 _05859_ vssd1 vssd1 vccd1 vccd1 _05860_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11077_ _04249_ net252 _04990_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12667__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14060__RESET_B net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _04342_ _04836_ _04946_ net263 vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__o211a_1
XANTENNA__08001__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10142__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12458__S net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11979_ _06181_ net292 net407 net2306 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11642__A1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ clknet_leaf_130_clk _00949_ net1176 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[706\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10445__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07941__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ clknet_leaf_105_clk _00880_ net1207 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[637\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07170_ final_design.cpu.reg_window\[650\] final_design.cpu.reg_window\[682\] net919
+ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08497__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11598__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12193__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_120_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07287__S net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12995__RESET_B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 _06125_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_4
Xfanout317 net318 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_8
X_09811_ _03259_ net443 net439 _03261_ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__o221a_1
Xfanout328 net330 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_8
Xfanout339 net342 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10381__B2 final_design.data_from_mem\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ _03198_ _03571_ _04495_ _03231_ net322 vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a221oi_1
X_06954_ final_design.cpu.reg_window\[529\] final_design.cpu.reg_window\[561\] net910
+ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__mux2_1
XANTENNA__07316__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _02837_ _04352_ _04591_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a21oi_1
X_06885_ _01832_ _01833_ _01834_ _01835_ net775 net796 vssd1 vssd1 vccd1 vccd1 _01836_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11330__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout274_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08624_ _03262_ _03574_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__nor2_1
XANTENNA__11780__B _05869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ net720 _03505_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__or2_1
XANTENNA__12368__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout441_A _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__A2 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout539_A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ _01911_ _02456_ _01912_ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08486_ net728 _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__or2_1
XANTENNA__13712__RESET_B net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08147__A _02030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10396__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07437_ net770 _02387_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout706_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout327_X net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1069_X net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07986__A _01939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08581__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07368_ final_design.cpu.reg_window\[707\] final_design.cpu.reg_window\[739\] net942
+ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09107_ _03715_ _03717_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__xor2_1
XANTENNA__11936__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06499__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07299_ final_design.cpu.reg_window\[261\] final_design.cpu.reg_window\[293\] net905
+ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_111_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_131_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09038_ _03788_ _03967_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold360 final_design.cpu.reg_window\[154\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 final_design.uart.BAUD_counter\[19\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 final_design.cpu.reg_window\[724\] vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net978 _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__nand2_1
XANTENNA__12361__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07925__S net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold393 final_design.cpu.reg_window\[366\] vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09762__B1 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__B2 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11447__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 net855 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_2
Xfanout851 net855 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_2
Xfanout862 net863 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_4
Xfanout873 net875 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_2
Xfanout884 net885 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09514__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07226__A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout895 _01437_ vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_4
X_12951_ clknet_leaf_55_clk _00189_ net1160 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_4
XANTENNA__11321__B1 _06014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1060 final_design.reqhand.instruction\[19\] vssd1 vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_172_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14120__Q final_design.VGA_data_control.v_count\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1071 final_design.cpu.reg_window\[623\] vssd1 vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902_ net204 net1890 net274 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__mux2_1
Xhold1082 final_design.cpu.reg_window\[276\] vssd1 vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12882_ clknet_leaf_87_clk _00120_ net1236 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[16\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold1093 final_design.cpu.reg_window\[868\] vssd1 vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ net195 net1959 net266 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__mux2_1
XANTENNA__10587__A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12416__A3 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11764_ net182 net2228 net418 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13503_ clknet_leaf_136_clk _00734_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[491\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07923__S0 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ net972 _05451_ _05453_ net968 vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11695_ net211 net635 vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__and2_1
X_13434_ clknet_leaf_150_clk _00665_ net1110 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[422\]
+ sky130_fd_sc_hd__dfrtp_1
X_10646_ _04767_ net254 vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__nor2_1
XANTENNA__08491__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11927__A2 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_102_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13365_ clknet_leaf_24_clk _00596_ net1158 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[353\]
+ sky130_fd_sc_hd__dfrtp_1
X_10577_ net813 _05320_ _05322_ net975 vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ net1843 net200 net364 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13296_ clknet_leaf_113_clk _00527_ net1212 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[284\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12247_ net594 _06176_ net504 _06273_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__a31o_1
XANTENNA__06799__X _01750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08100__S0 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__A2 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11865__B net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ net2094 net207 net381 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__mux2_1
XANTENNA__10363__B2 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14140__1257 vssd1 vssd1 vccd1 vccd1 _14140__1257/HI net1257 sky130_fd_sc_hd__conb_1
X_11129_ net816 _05839_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_25 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_169_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_169_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_161_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06670_ final_design.cpu.reg_window\[538\] final_design.cpu.reg_window\[570\] net952
+ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__mux2_1
XANTENNA__12188__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08340_ net538 _03289_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__or2_1
XANTENNA__10418__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08271_ _03218_ _03219_ _03220_ _03221_ net686 net700 vssd1 vssd1 vccd1 vccd1 _03222_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11820__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07222_ final_design.cpu.reg_window\[648\] final_design.cpu.reg_window\[680\] net920
+ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06914__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07047__A1 final_design.data_from_mem\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07153_ final_design.cpu.reg_window\[330\] final_design.cpu.reg_window\[362\] net921
+ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ final_design.cpu.reg_window\[268\] final_design.cpu.reg_window\[300\] net927
+ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__A0 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12343__A2 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06502__X _01453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout391_A _06265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__B2 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06869__B _01468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11551__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07986_ _01939_ net617 vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_35_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09725_ net555 net554 net553 net552 net454 net463 vssd1 vssd1 vccd1 vccd1 _04644_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10106__A1 final_design.VGA_data_control.v_count\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_06937_ final_design.cpu.reg_window\[273\] final_design.cpu.reg_window\[305\] net918
+ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__mux2_1
XANTENNA__11303__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout656_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09656_ net80 _04189_ net81 vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__o21ai_1
X_06868_ net751 net854 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__nand2_1
XANTENNA__08576__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09261__A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _03555_ _03556_ _03488_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a21o_1
XANTENNA__12098__S net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout823_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _03164_ _04505_ _03162_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__a21oi_1
X_06799_ net894 _01731_ _01737_ _01743_ _01749_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__o32a_4
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10409__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08538_ final_design.cpu.reg_window\[321\] final_design.cpu.reg_window\[353\] net854
+ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07905__S0 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08469_ net625 _03415_ _03416_ net533 vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_147_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10500_ _05233_ _05246_ _05244_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__o21bai_2
XTAP_TAPCELL_ROW_133_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09027__A2 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11480_ _06017_ net2463 net309 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08605__A _02390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10431_ _03613_ _05180_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__or2_2
XFILLER_0_123_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12031__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire559 _01626_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_150_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12127__A _06094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07133__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13150_ clknet_leaf_21_clk _00381_ net1124 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[138\]
+ sky130_fd_sc_hd__dfrtp_1
X_10362_ net4 net1036 net1019 final_design.data_from_mem\[11\] vssd1 vssd1 vccd1 vccd1
+ _00115_ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14115__Q final_design.reqhand.data_from_UART\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12101_ net2067 net237 net388 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__mux2_1
XANTENNA__11790__B1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ net1061 _05146_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__nand2_1
X_13081_ clknet_leaf_167_clk _00312_ net1081 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12334__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ net2004 net223 net396 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__mux2_1
Xhold190 final_design.VGA_data_control.ready_data\[10\] vssd1 vssd1 vccd1 vccd1 net1543
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11685__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08340__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__B2 final_design.data_from_mem\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10896__A2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout670 _02511_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_4
Xfanout681 _02328_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_2
Xfanout692 net698 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_4
X_13983_ clknet_leaf_135_clk _01214_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[971\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11905__S net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ clknet_leaf_33_clk _00172_ net1129 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13634__RESET_B net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07390__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12865_ clknet_leaf_82_clk _00103_ net1248 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11206__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ net224 net2362 net266 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12270__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11747_ net214 net2461 net418 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07372__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06734__S net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11678_ net585 net423 _06197_ net297 net1640 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__a32o_1
XFILLER_0_126_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13417_ clknet_leaf_89_clk _00648_ net1231 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[405\]
+ sky130_fd_sc_hd__dfrtp_1
X_10629_ net98 final_design.VGA_adr\[6\] _05370_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10033__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ clknet_leaf_100_clk _00579_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[336\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13279_ clknet_leaf_137_clk _00510_ net1169 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[267\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09726__A0 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07565__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09346__A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__B2 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ final_design.cpu.reg_window\[725\] final_design.cpu.reg_window\[757\] net885
+ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07752__A2 _02698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12089__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ final_design.cpu.reg_window\[984\] final_design.cpu.reg_window\[1016\] net869
+ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11815__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ _04427_ _04428_ net448 vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__a21o_1
X_06722_ _01669_ _01670_ _01671_ _01672_ net785 net803 vssd1 vssd1 vccd1 vccd1 _01673_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_91_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06909__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10939__B _05662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06938__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09441_ _02738_ _03594_ _04359_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__a21o_1
X_06653_ final_design.cpu.reg_window\[474\] final_design.cpu.reg_window\[506\] net955
+ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09372_ _02609_ _04050_ _03605_ _02573_ _02575_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06584_ net900 _01528_ _01534_ _01521_ _01522_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__a32oi_1
XFILLER_0_86_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08323_ net727 _03273_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout237_A _05904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08560__S0 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08254_ _03201_ _03202_ _03203_ _03204_ net690 net710 vssd1 vssd1 vccd1 vccd1 _03205_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07205_ net896 _02148_ _02154_ _02141_ _02142_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a32o_1
XFILLER_0_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08185_ final_design.cpu.reg_window\[334\] final_design.cpu.reg_window\[366\] net852
+ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout404_A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10024__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07136_ final_design.cpu.reg_window\[587\] final_design.cpu.reg_window\[619\] net937
+ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07067_ final_design.cpu.reg_window\[653\] final_design.cpu.reg_window\[685\] net915
+ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__mux2_1
XANTENNA__12381__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10327__B2 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A _01426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08940__A1 final_design.CPU_instr_adr\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ final_design.cpu.reg_window\[849\] final_design.cpu.reg_window\[881\] net836
+ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _03070_ _04504_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__nand2_1
X_10980_ net975 _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09639_ _02997_ net446 net442 _02994_ _04557_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__o221a_2
XFILLER_0_167_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12650_ _06312_ net1484 net994 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11601_ net580 net422 _06156_ net304 net1702 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__a32o_1
XANTENNA__11055__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12252__A1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12581_ _01395_ net1014 vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__nor2_2
XANTENNA__10865__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07354__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11532_ net1725 net183 net526 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14251_ net1316 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XANTENNA__08208__B1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11463_ net217 net2412 net308 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13202_ clknet_leaf_38_clk _00433_ net1135 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[190\]
+ sky130_fd_sc_hd__dfrtp_1
X_10414_ _05176_ _05180_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__or2_4
XANTENNA__11212__C1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12555__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__B1 _04124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14182_ clknet_leaf_56_clk _01356_ net1163 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11394_ _01507_ net650 _06078_ net653 vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13133_ clknet_leaf_103_clk _00364_ net1201 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10345_ net1493 net1024 net1001 final_design.data_from_mem\[30\] vssd1 vssd1 vccd1
+ vccd1 _00102_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07385__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__A2 _02929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13064_ clknet_leaf_126_clk _00295_ net1192 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_10276_ final_design.uart.BAUD_counter\[28\] _05134_ net812 vssd1 vssd1 vccd1 vccd1
+ _05136_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10318__B2 final_design.data_from_mem\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07719__C1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12015_ _06217_ net284 net401 net1922 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__a22o_1
XANTENNA__09723__A3 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13815__RESET_B net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11279__C1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13966_ clknet_leaf_114_clk _01197_ net1210 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[954\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06729__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09105__S net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12917_ clknet_leaf_33_clk _00155_ net1129 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07042__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13897_ clknet_leaf_88_clk _01128_ net1237 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[885\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12848_ clknet_leaf_78_clk _00086_ net1250 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08944__S net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12243__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08542__S0 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12546__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold904 final_design.cpu.reg_window\[644\] vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold915 final_design.cpu.reg_window\[483\] vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 final_design.cpu.reg_window\[743\] vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold937 final_design.cpu.reg_window\[866\] vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 final_design.cpu.reg_window\[805\] vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10714__S net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold959 final_design.cpu.reg_window\[894\] vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ _02736_ net444 vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06856__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08941_ _03762_ _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08872_ _03801_ _03820_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__or2_1
XANTENNA__06987__X _01938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07823_ final_design.cpu.reg_window\[213\] final_design.cpu.reg_window\[245\] net884
+ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__mux2_1
XANTENNA__07281__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout187_A _06052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11772__C net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07754_ _02704_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__inv_2
XANTENNA__06639__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06705_ net771 _01655_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07685_ _01507_ net626 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout354_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09424_ net492 _04205_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06636_ final_design.cpu.reg_window\[923\] final_design.cpu.reg_window\[955\] net961
+ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12234__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ _04074_ _04264_ _04273_ _04263_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__o211a_1
XANTENNA__12376__S net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06567_ final_design.cpu.reg_window\[221\] final_design.cpu.reg_window\[253\] net959
+ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout521_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout619_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08989__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07336__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ net889 _03238_ _03244_ _03250_ _03256_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__o32a_4
X_09286_ net482 _04204_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__or2_2
X_06498_ final_design.cpu.reg_window\[542\] final_design.cpu.reg_window\[574\] net931
+ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08237_ final_design.cpu.reg_window\[587\] final_design.cpu.reg_window\[619\] net857
+ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08168_ final_design.cpu.reg_window\[783\] final_design.cpu.reg_window\[815\] net824
+ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout890_A _01687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11745__A0 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07119_ final_design.cpu.reg_window\[459\] final_design.cpu.reg_window\[491\] net938
+ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08099_ final_design.cpu.reg_window\[140\] final_design.cpu.reg_window\[172\] net847
+ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10130_ _05002_ _05035_ final_design.v_out vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_state\[0\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10061_ _04325_ _04326_ _04964_ _04966_ _04979_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_73_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07177__A0 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07933__S net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__C1 _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13226__RESET_B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout943_X net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__S net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13820_ clknet_leaf_144_clk _01051_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[808\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_162_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13751_ clknet_leaf_143_clk _00982_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[739\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07024__S0 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ net52 _05688_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_82_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12702_ final_design.VGA_data_control.v_count\[5\] _06337_ _06342_ vssd1 vssd1 vccd1
+ vccd1 _06343_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_97_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10484__B1 _04990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07575__S1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13682_ clknet_leaf_41_clk _00913_ net1150 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[670\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10894_ _05600_ _05621_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12633_ final_design.VGA_data_control.ready_data\[4\] net1035 net990 final_design.data_from_mem\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08336__Y _03287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12564_ net1065 final_design.uart.working_data\[2\] vssd1 vssd1 vccd1 vccd1 _06287_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_93_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11984__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11515_ net2241 net209 net524 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__mux2_1
X_12495_ _06155_ net350 net332 net2212 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14234_ net1299 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_151_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12528__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ net228 net646 vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14165_ clknet_leaf_78_clk _01339_ net1250 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08601__B1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11377_ final_design.data_from_mem\[28\] net235 net233 vssd1 vssd1 vccd1 vccd1 _06064_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13116_ clknet_leaf_148_clk _00347_ net1126 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_10328_ net1523 net1022 net999 final_design.data_from_mem\[13\] vssd1 vssd1 vccd1
+ vccd1 _00085_ sky130_fd_sc_hd__a22o_1
X_14096_ clknet_leaf_84_clk _01293_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09157__A1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13047_ clknet_leaf_144_clk _00278_ net1182 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_10259_ _05124_ _05125_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__nor2_1
Xfanout1240 net1243 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07843__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1251 net1255 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09624__A _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08117__C1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13949_ clknet_leaf_12_clk _01180_ net1093 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[937\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_73_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12949__RESET_B net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10475__B1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07470_ _01480_ net738 _02095_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06421_ final_design.reqhand.instruction\[4\] vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09140_ _04057_ _04058_ net479 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__mux2_1
XANTENNA__09093__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11975__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_62_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09071_ net2555 net1028 _03997_ vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12519__A2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08022_ final_design.cpu.reg_window\[83\] final_design.cpu.reg_window\[115\] net825
+ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold701 final_design.cpu.reg_window\[942\] vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold712 final_design.cpu.reg_window\[1009\] vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold723 final_design.cpu.reg_window\[667\] vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold734 final_design.cpu.reg_window\[959\] vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 final_design.cpu.reg_window\[554\] vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 final_design.cpu.reg_window\[171\] vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A2 _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold767 final_design.cpu.reg_window\[393\] vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 final_design.cpu.reg_window\[406\] vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09973_ net483 _04891_ _04341_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold789 final_design.cpu.reg_window\[675\] vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09148__A1 _04066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ net629 _03864_ _03866_ net258 vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout1011_A _06295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09699__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08855_ _03783_ _03805_ final_design.CPU_instr_adr\[31\] net1049 vssd1 vssd1 vccd1
+ vccd1 _00242_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout471_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07806_ final_design.cpu.reg_window\[729\] final_design.cpu.reg_window\[761\] net859
+ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08786_ _03734_ _03736_ _03686_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11258__A2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07737_ final_design.cpu.reg_window\[794\] final_design.cpu.reg_window\[826\] net872
+ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__mux2_1
XANTENNA__12455__A1 net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout736_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__B1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07668_ final_design.cpu.reg_window\[222\] final_design.cpu.reg_window\[254\] net848
+ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07331__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09407_ net89 _04195_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__xor2_1
X_06619_ _01477_ _01497_ net672 _01569_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a211o_2
XANTENNA__12207__A1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07882__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout903_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07599_ final_design.cpu.reg_window\[285\] final_design.cpu.reg_window\[317\] net880
+ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09338_ net622 _03549_ _03523_ _01453_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__a211o_1
XFILLER_0_106_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11966__B1 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09269_ net76 net77 _04187_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__or3_1
XANTENNA__10604__A_N net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11300_ net654 net202 vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__and2_1
XANTENNA__07928__S net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12280_ net594 _06210_ net518 net371 net1834 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__a32o_1
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11718__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout893_X net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11231_ net582 net422 _05935_ net316 net1965 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_75_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11162_ _04879_ _05143_ net600 _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_112_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09139__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ net1064 _05023_ _05003_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__o21ai_1
X_11093_ _05813_ _05814_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_164_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07663__S net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _04249_ _04252_ _04289_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__a21boi_1
XANTENNA__11693__B net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 final_design.VGA_data_control.data_to_VGA\[29\] vssd1 vssd1 vccd1 vccd1 net1403
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 final_design.reqhand.data_from_UART\[6\] vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold72 final_design.reqhand.instruction\[30\] vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 net141 vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 final_design.VGA_data_control.data_to_VGA\[5\] vssd1 vssd1 vccd1 vccd1 net1447
+ sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ clknet_leaf_18_clk _01034_ net1121 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[791\]
+ sky130_fd_sc_hd__dfrtp_1
X_11995_ _06197_ net289 net402 net2268 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_55_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11913__S net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13734_ clknet_leaf_171_clk _00965_ net1075 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[722\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07899__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10946_ _04918_ net254 vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__nor2_1
XANTENNA__08494__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_119_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13665_ clknet_leaf_159_clk _00896_ net1106 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[653\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10472__A3 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ _04598_ net254 vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11214__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ final_design.uart.working_data\[3\] net1401 _05080_ vssd1 vssd1 vccd1 vccd1
+ _01309_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ clknet_leaf_152_clk _00827_ net1116 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[584\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10304__S0 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12547_ _06210_ net358 net326 net2159 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07838__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12478_ _06138_ net347 net331 net1857 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14217_ net1286 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
X_11429_ net2202 net199 net311 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__mux2_1
XANTENNA__09378__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13830__RESET_B net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08242__B net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14148_ clknet_leaf_82_clk _01322_ net1247 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14079_ clknet_leaf_72_clk _01276_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_06970_ final_design.cpu.reg_window\[144\] final_design.cpu.reg_window\[176\] net958
+ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__mux2_1
XANTENNA__12134__A0 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07573__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12685__B2 final_design.data_from_mem\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1070 net1071 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_4
Xfanout1081 net1083 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_4
X_08640_ _02932_ _02933_ _03586_ _03588_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__o22a_1
XFILLER_0_174_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1092 net1094 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__clkbuf_4
X_08571_ _03520_ _03521_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_46_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11823__S net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07522_ _01631_ _02471_ _01600_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10999__A1 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10999__B2 _04040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07453_ final_design.cpu.reg_window\[128\] final_design.cpu.reg_window\[160\] net943
+ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__mux2_1
XANTENNA__11660__A2 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06404_ final_design.CPU_instr_adr\[27\] vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
XANTENNA__11124__A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07384_ final_design.cpu.reg_window\[450\] final_design.cpu.reg_window\[482\] net947
+ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11948__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13989__RESET_B net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09123_ net1007 net1003 vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__nor2_4
XFILLER_0_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08704__Y _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout317_A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1059_A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09054_ _03980_ _03982_ final_design.CPU_instr_adr\[9\] net1049 vssd1 vssd1 vccd1
+ vccd1 _00220_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06652__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12951__Q net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08005_ final_design.cpu.reg_window\[656\] final_design.cpu.reg_window\[688\] net879
+ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__mux2_1
XANTENNA__11130__Y _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold520 final_design.uart.working_data\[5\] vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 final_design.cpu.reg_window\[548\] vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold542 final_design.cpu.reg_window\[374\] vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1226_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold553 final_design.cpu.reg_window\[863\] vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold564 final_design.cpu.reg_window\[253\] vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 final_design.cpu.reg_window\[918\] vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold586 final_design.cpu.reg_window\[497\] vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 final_design.cpu.reg_window\[69\] vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11794__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09956_ _03488_ _03555_ _03556_ _04124_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08579__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1014_X net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08907_ final_design.CPU_instr_adr\[24\] _03797_ final_design.CPU_instr_adr\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__a21oi_1
X_09887_ net733 _04805_ net79 vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__o21ai_1
Xhold1220 final_design.vga.v_current_state\[1\] vssd1 vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ final_design.CPU_instr_adr\[11\] _03788_ vssd1 vssd1 vccd1 vccd1 _03789_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07778__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ _03710_ _03719_ _03709_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__a21o_1
XFILLER_0_169_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10800_ final_design.CPU_instr_adr\[17\] _05534_ net1066 vssd1 vssd1 vccd1 vccd1
+ _05535_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06827__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11780_ net656 _05869_ net220 vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_68_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08608__A _02356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10731_ _05464_ _05468_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11034__A _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13450_ clknet_leaf_2_clk _00681_ net1079 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[438\]
+ sky130_fd_sc_hd__dfrtp_1
X_10662_ _05347_ _05385_ _05403_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11939__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12401_ _06099_ net353 net341 net2446 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07607__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13381_ clknet_leaf_149_clk _00612_ net1119 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[369\]
+ sky130_fd_sc_hd__dfrtp_1
X_10593_ _05336_ _05337_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__nor2_1
XANTENNA__12600__B2 final_design.data_from_mem\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12332_ net2532 net361 net350 _05865_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06562__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12263_ net679 _06193_ _06262_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11167__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14002_ clknet_leaf_26_clk _01233_ net1142 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[990\]
+ sky130_fd_sc_hd__dfrtp_1
X_11214_ net598 _05919_ _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__and3_1
X_12194_ net2173 net179 net381 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__mux2_1
XANTENNA__07466__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ net670 _04028_ net746 vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08489__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09174__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_X net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07218__S0 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ _05757_ _05775_ _05792_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__o31ai_2
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12667__B2 final_design.data_from_mem\[21\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ _02837_ net446 _04943_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_127_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_28_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11978_ _06180_ net290 net406 net1979 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10929_ net1069 _05656_ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__a21oi_1
X_13717_ clknet_leaf_25_clk _00948_ net1144 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[705\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_152_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07141__B net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07941__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13648_ clknet_leaf_104_clk _00879_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[636\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12198__A3 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13579_ clknet_leaf_15_clk _00810_ net1102 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[567\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10602__B1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_167_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07568__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11598__B net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11158__A1 net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12355__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10007__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11818__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout307 net310 vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_6
X_09810_ _03262_ _04087_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__nand2_1
Xfanout318 _05851_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06585__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout329 net330 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_8
X_09741_ _03230_ _04495_ _03571_ _03198_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a211o_1
X_06953_ final_design.cpu.reg_window\[593\] final_design.cpu.reg_window\[625\] net910
+ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07316__B _01659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _02803_ _03034_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__nand2_1
XANTENNA__10023__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06884_ final_design.cpu.reg_window\[147\] final_design.cpu.reg_window\[179\] net908
+ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_145_Left_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08623_ _02185_ _03289_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__nand2_1
XANTENNA__10958__A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11881__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout267_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ _03501_ _03502_ _03503_ _03504_ net687 net708 vssd1 vssd1 vccd1 vccd1 _03505_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07505_ _01941_ _02455_ _01940_ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a21oi_1
X_08485_ _03432_ _03433_ _03434_ _03435_ net692 net711 vssd1 vssd1 vccd1 vccd1 _03436_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout434_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10396__C net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07436_ _02383_ _02384_ _02385_ _02386_ net781 net792 vssd1 vssd1 vccd1 vccd1 _02387_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07051__B _02000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10693__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07986__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12384__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07367_ net764 _02317_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout601_A _05199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09106_ net1031 _04027_ net1050 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__mux2_1
XANTENNA__09259__A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06499__S1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07298_ final_design.cpu.reg_window\[325\] final_design.cpu.reg_window\[357\] net905
+ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09037_ final_design.CPU_instr_adr\[9\] _03787_ final_design.CPU_instr_adr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_131_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12775__6 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__inv_2
XFILLER_0_13_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12346__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1229_X net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08014__A1 _01908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold350 final_design.cpu.reg_window\[850\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 final_design.cpu.reg_window\[178\] vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 final_design.cpu.reg_window\[156\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 net132 vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold394 final_design.cpu.reg_window\[640\] vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout830 net835 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08970__C1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout841 net842 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_4
Xfanout852 net853 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_4
X_09939_ net264 _04854_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__and3_1
XANTENNA__12649__B2 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 net864 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_4
Xfanout874 net875 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_4
Xfanout885 net886 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__clkbuf_2
X_12950_ clknet_leaf_55_clk _00188_ net1160 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_1
Xfanout896 net897 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_8
Xhold1050 final_design.cpu.reg_window\[67\] vssd1 vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 final_design.cpu.reg_window\[1021\] vssd1 vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net221 net1936 net276 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__mux2_1
Xhold1072 final_design.cpu.reg_window\[418\] vssd1 vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ clknet_leaf_79_clk _00119_ net1249 vssd1 vssd1 vccd1 vccd1 final_design.data_from_mem\[15\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold1083 final_design.cpu.reg_window\[705\] vssd1 vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10868__A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1094 final_design.cpu.reg_window\[290\] vssd1 vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11463__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _06017_ net2294 net269 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10587__B final_design.VGA_adr\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07242__A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11763_ net185 net1974 net419 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__mux2_1
XANTENNA__11624__A2 net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10832__B1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10714_ final_design.CPU_instr_adr\[13\] _03951_ net1070 vssd1 vssd1 vccd1 vccd1
+ _05453_ sky130_fd_sc_hd__mux2_1
XANTENNA__07923__S1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13502_ clknet_leaf_22_clk _00733_ net1123 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[490\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11694_ net432 net583 _06205_ net297 net1896 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13433_ clknet_leaf_165_clk _00664_ net1085 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[421\]
+ sky130_fd_sc_hd__dfrtp_1
X_10645_ net1015 _05384_ _05387_ net1042 net1736 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__a32o_1
XFILLER_0_119_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11388__A1 _04324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07388__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13364_ clknet_leaf_103_clk _00595_ net1186 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[352\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_691 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10576_ net971 _05319_ _05321_ net969 vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__o22a_1
XANTENNA__09450__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12315_ net2017 net202 net364 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13295_ clknet_leaf_91_clk _00526_ net1232 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[283\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12337__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12246_ final_design.cpu.reg_window\[720\] net375 vssd1 vssd1 vccd1 vccd1 _06273_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_139_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08100__S1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__Y _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ net1940 net210 net380 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__mux2_1
XANTENNA__09616__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ net816 _05839_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__nor2_8
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08308__A2 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059_ _05780_ _05781_ _05761_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08947__S net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11312__A1 final_design.data_from_mem\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09632__A net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09351__B _04094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10823__B1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08270_ final_design.cpu.reg_window\[522\] final_design.cpu.reg_window\[554\] net837
+ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07221_ final_design.cpu.reg_window\[712\] final_design.cpu.reg_window\[744\] net921
+ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07152_ final_design.cpu.reg_window\[394\] final_design.cpu.reg_window\[426\] net936
+ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07083_ final_design.cpu.reg_window\[332\] final_design.cpu.reg_window\[364\] net929
+ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_160_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__A1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10354__A2 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11551__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07985_ _02935_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout384_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ _04641_ _04642_ net477 vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__mux2_1
X_06936_ final_design.cpu.reg_window\[337\] final_design.cpu.reg_window\[369\] net918
+ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__mux2_1
XANTENNA__11303__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09655_ _04571_ _04573_ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06867_ _01816_ _01817_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__nand2_1
XANTENNA__12379__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout551_A _01850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11854__A2 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout649_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _03555_ _03556_ _03488_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11136__X _05851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09261__B net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _03070_ _03101_ _04504_ _04137_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__a31o_1
Xclkbuf_3_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_clk sky130_fd_sc_hd__clkbuf_8
X_06798_ net758 _01748_ net894 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_65_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08537_ _03486_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__nor2_2
XANTENNA__10200__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07905__S1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07997__A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08468_ net625 _03415_ _03416_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__a21o_1
X_07419_ final_design.cpu.reg_window\[65\] final_design.cpu.reg_window\[97\] net931
+ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08399_ _03346_ _03347_ _03348_ _03349_ net685 net699 vssd1 vssd1 vccd1 vccd1 _03350_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_162_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08605__B _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10430_ net1478 net1040 _05198_ net247 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12127__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10361_ net3 net1038 net1021 final_design.data_from_mem\[10\] vssd1 vssd1 vccd1 vccd1
+ _00114_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12100_ net1869 net223 net388 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09717__A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13080_ clknet_leaf_133_clk _00311_ net1174 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06840__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10292_ _05144_ _05145_ _01384_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout973_X net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ net2184 net239 net398 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__mux2_1
Xhold180 final_design.cpu.reg_window\[190\] vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold191 net163 vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_109_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout660 _05143_ vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__buf_4
Xfanout682 net684 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_8
Xfanout693 net695 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_8
X_13982_ clknet_leaf_19_clk _01213_ net1120 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[970\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ clknet_leaf_34_clk _00171_ net1133 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ clknet_leaf_81_clk _00102_ net1247 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11815_ net240 net2429 net268 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__mux2_1
XANTENNA_output101_A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ net216 net1930 net417 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ net226 net636 vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12558__B1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11222__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10628_ _05351_ _05370_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13416_ clknet_leaf_117_clk _00647_ net1194 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[404\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12022__A2 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13347_ clknet_leaf_4_clk _00578_ net1086 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[335\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10559_ _05268_ _05305_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11781__B2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13278_ clknet_leaf_22_clk _00509_ net1127 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[266\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09726__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ net679 _06158_ _06262_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10336__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11533__A1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__A _02097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07832__S0 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ final_design.cpu.reg_window\[792\] final_design.cpu.reg_window\[824\] net869
+ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06721_ final_design.cpu.reg_window\[408\] final_design.cpu.reg_window\[440\] net949
+ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09440_ _02769_ _03597_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__nand2_1
X_06652_ final_design.cpu.reg_window\[282\] final_design.cpu.reg_window\[314\] net955
+ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09371_ _04286_ _04288_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_82_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06583_ net773 _01533_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11831__S net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ _03269_ _03270_ _03271_ _03272_ net686 net707 vssd1 vssd1 vccd1 vccd1 _03273_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06925__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08253_ final_design.cpu.reg_window\[394\] final_design.cpu.reg_window\[426\] net854
+ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__mux2_1
XANTENNA__08560__S1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12549__B1 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07204_ net896 _02148_ _02154_ _02141_ _02142_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12013__A2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08184_ _02000_ net604 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__nand2_1
XANTENNA__09414__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07135_ final_design.cpu.reg_window\[651\] final_design.cpu.reg_window\[683\] net938
+ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10971__A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1041_A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1139_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07066_ final_design.cpu.reg_window\[717\] final_design.cpu.reg_window\[749\] net915
+ vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07440__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10035__X _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10327__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07057__A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ final_design.cpu.reg_window\[913\] final_design.cpu.reg_window\[945\] net836
+ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__mux2_1
XANTENNA__08587__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06919_ final_design.cpu.reg_window\[786\] final_design.cpu.reg_window\[818\] net901
+ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__mux2_1
X_09707_ _04124_ _04625_ _04624_ net263 vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout933_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07899_ net726 _02849_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09638_ _02995_ net441 vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__nand2_1
XANTENNA__07900__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ net320 _04487_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11741__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ net177 net643 vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__and2_1
XFILLER_0_167_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12580_ _01395_ _04037_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11531_ net1709 net184 net527 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14250_ net1315 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11462_ net218 net648 vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__and2_1
XANTENNA__08208__A1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12004__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13201_ clknet_leaf_107_clk _00432_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[189\]
+ sky130_fd_sc_hd__dfrtp_1
X_10413_ net1544 net1040 _05189_ net247 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__a22o_1
X_14181_ clknet_leaf_68_clk _01355_ net1222 vssd1 vssd1 vccd1 vccd1 final_design.VGA_adr\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11393_ final_design.data_from_mem\[30\] net236 net234 vssd1 vssd1 vccd1 vccd1 _06078_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13132_ clknet_leaf_122_clk _00363_ net1197 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input62_A mem_adr_start[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ net1475 net1023 net1000 final_design.data_from_mem\[29\] vssd1 vssd1 vccd1
+ vccd1 _00101_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_78_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13063_ clknet_leaf_8_clk _00294_ net1087 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10275_ _05134_ _05135_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__nor2_1
X_12014_ _06216_ net278 net400 net1982 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_167_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11916__S net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10820__S net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout490 net492 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11279__B1 _05976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13965_ clknet_leaf_128_clk _01196_ net1180 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[953\]
+ sky130_fd_sc_hd__dfrtp_1
X_12916_ clknet_leaf_159_clk _00154_ net1106 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07042__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ clknet_leaf_119_clk _01127_ net1200 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[884\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12491__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09892__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12847_ clknet_leaf_78_clk _00085_ net1247 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.ready_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12798__29 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__inv_2
XFILLER_0_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08542__S1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11729_ net180 net637 vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09086__A1_N net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold905 final_design.cpu.reg_window\[167\] vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold916 final_design.cpu.reg_window\[501\] vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 final_design.cpu.reg_window\[806\] vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06480__S net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold938 final_design.cpu.reg_window\[1011\] vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 final_design.cpu.reg_window\[114\] vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06856__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08940_ final_design.CPU_instr_adr\[20\] _01823_ _03753_ vssd1 vssd1 vccd1 vccd1
+ _03881_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11506__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08871_ final_design.CPU_instr_adr\[29\] _03800_ vssd1 vssd1 vccd1 vccd1 _03820_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07805__S0 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11826__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07822_ _01788_ net608 vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07281__S1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07753_ _02701_ _02703_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__nor2_1
XANTENNA__11809__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06704_ _01651_ _01652_ _01653_ _01654_ net783 net793 vssd1 vssd1 vccd1 vccd1 _01655_
+ sky130_fd_sc_hd__mux4_1
X_07684_ _02622_ _02623_ _02634_ net889 vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12482__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09423_ net603 _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__or2_4
X_06635_ final_design.cpu.reg_window\[987\] final_design.cpu.reg_window\[1019\] net961
+ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__mux2_1
XANTENNA__11690__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__A _05673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout347_A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09354_ net492 _04231_ _04261_ _04265_ _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__o311a_1
XFILLER_0_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06566_ final_design.cpu.reg_window\[29\] final_design.cpu.reg_window\[61\] net959
+ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08305_ net719 _03255_ net889 vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07379__A2_N net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09285_ net530 net459 _04203_ net469 vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06497_ final_design.cpu.reg_window\[606\] final_design.cpu.reg_window\[638\] net931
+ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout514_A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1256_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ final_design.cpu.reg_window\[651\] final_design.cpu.reg_window\[683\] net857
+ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08167_ final_design.cpu.reg_window\[847\] final_design.cpu.reg_window\[879\] net827
+ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__mux2_1
XANTENNA__12392__S net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_X net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09267__A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ final_design.cpu.reg_window\[267\] final_design.cpu.reg_window\[299\] net938
+ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08098_ final_design.cpu.reg_window\[204\] final_design.cpu.reg_window\[236\] net846
+ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout883_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07049_ net750 net673 _01851_ _01999_ _01821_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10060_ _04967_ _04969_ _04977_ _04978_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_73_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07177__A1 _01505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12170__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11736__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout936_X net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11037__A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ _05689_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__inv_2
X_13750_ clknet_leaf_130_clk _00981_ net1190 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[738\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12473__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07024__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12701_ final_design.VGA_data_control.v_count\[5\] _06339_ _06335_ vssd1 vssd1 vccd1
+ vccd1 _06342_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10484__A1 _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09730__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10893_ _05606_ _05622_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__or2_1
X_13681_ clknet_leaf_106_clk _00912_ net1208 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[669\]
+ sky130_fd_sc_hd__dfrtp_1
X_12632_ _06303_ net1517 net992 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12563_ net1065 _05078_ _05066_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11514_ net1636 net211 net525 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09729__X _04648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12494_ _06154_ net358 net334 net1860 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14233_ net1298 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11445_ net232 net2378 net310 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07396__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14164_ clknet_leaf_81_clk _01338_ net1247 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11376_ net740 _03829_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ net1481 net1023 net1000 final_design.data_from_mem\[12\] vssd1 vssd1 vccd1
+ vccd1 _00084_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ clknet_leaf_156_clk _00346_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_14095_ clknet_leaf_84_clk _01292_ net1228 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13046_ clknet_leaf_130_clk _00277_ net1175 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09157__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10258_ net2574 _05123_ net809 vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_147_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1230 net1231 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_4
Xfanout1241 net1242 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1252 net1253 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__clkbuf_4
X_10189_ _05078_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__inv_2
XANTENNA__12331__A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13948_ clknet_leaf_148_clk _01179_ net1125 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[936\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06679__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10475__B2 final_design.CPU_instr_adr\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10786__A net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13879_ clknet_leaf_141_clk _01110_ net1184 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[867\]
+ sky130_fd_sc_hd__dfrtp_1
X_06420_ final_design.data_from_mem\[2\] vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12989__RESET_B net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09093__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09070_ _03655_ _03995_ _03996_ _03993_ net1049 vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__o221a_1
XANTENNA__09639__X _04558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08021_ net718 _02971_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold702 final_design.cpu.reg_window\[506\] vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold713 final_design.cpu.reg_window\[873\] vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_1__f_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold724 final_design.cpu.reg_window\[947\] vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold735 final_design.cpu.reg_window\[936\] vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 final_design.cpu.reg_window\[445\] vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 final_design.cpu.reg_window\[769\] vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 final_design.cpu.reg_window\[39\] vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold779 final_design.cpu.reg_window\[884\] vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _04663_ _04815_ net471 vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08923_ net629 _03865_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13777__RESET_B net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11409__X _06092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout297_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__A3 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10313__X _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ net260 _03804_ net1029 vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07805_ _02752_ _02753_ _02754_ _02755_ net693 net712 vssd1 vssd1 vccd1 vccd1 _02756_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11128__Y _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08785_ _01365_ _02063_ _03685_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ final_design.cpu.reg_window\[858\] final_design.cpu.reg_window\[890\] net872
+ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08659__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09550__A _04072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__B2 final_design.CPU_instr_adr\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ final_design.cpu.reg_window\[30\] final_design.cpu.reg_window\[62\] net847
+ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12387__S net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout252_X net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout631_A _02506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__A1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout729_A _01720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09406_ net734 _04324_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__nor2_2
XFILLER_0_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06618_ net753 _01568_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07882__A2 _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07598_ final_design.cpu.reg_window\[349\] final_design.cpu.reg_window\[381\] net880
+ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06549_ final_design.reqhand.instruction\[31\] net983 vssd1 vssd1 vccd1 vccd1 _01500_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_35_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09337_ _03602_ _04254_ _02673_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout1161_X net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ net75 _04186_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08219_ final_design.cpu.reg_window\[267\] final_design.cpu.reg_window\[299\] net857
+ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10635__S net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09199_ net491 net319 vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11718__A1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11179__C1 _05889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ net655 net215 vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__and2_2
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08044__C1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08105__S net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11161_ net665 _05871_ _05873_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10112_ _05023_ _05024_ _05006_ vssd1 vssd1 vccd1 vccd1 final_design.vga.v_next_count\[3\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__09139__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11092_ net59 _05799_ _05810_ _05812_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_164_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11466__S net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ _04571_ _04573_ _04388_ _04425_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__o211a_1
Xhold40 final_design.VGA_data_control.data_to_VGA\[14\] vssd1 vssd1 vccd1 vccd1 net1393
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 final_design.cpu.reg_window\[4\] vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _01313_ vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold73 final_design.cpu.reg_window\[735\] vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 final_design.reqhand.instruction\[24\] vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 final_design.cpu.reg_window\[200\] vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ clknet_leaf_164_clk _01033_ net1084 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[790\]
+ sky130_fd_sc_hd__dfrtp_1
X_11994_ net2520 net402 _06258_ net434 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__a22o_1
XANTENNA__11654__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13733_ clknet_leaf_4_clk _00964_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[721\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10457__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10945_ _05508_ _05672_ _05671_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__o21bai_4
XANTENNA__12297__S net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13664_ clknet_leaf_44_clk _00895_ net1146 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[652\]
+ sky130_fd_sc_hd__dfrtp_1
X_10876_ net1015 _05606_ _05607_ net1043 net1467 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12615_ net1406 final_design.reqhand.data_from_UART\[1\] _05080_ vssd1 vssd1 vccd1
+ vccd1 _01308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13595_ clknet_leaf_156_clk _00826_ net1114 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[583\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10304__S1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12546_ _06209_ net345 net323 net2200 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12477_ _06137_ net349 net332 net1985 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11230__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_4 _02961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ net1285 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
X_11428_ net1881 net201 net311 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14147_ clknet_leaf_72_clk _01321_ net1247 vssd1 vssd1 vccd1 vccd1 final_design.VGA_data_control.data_to_VGA\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11359_ net748 _03844_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09906__Y _04825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10393__B1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14078_ clknet_leaf_72_clk _01275_ net1241 vssd1 vssd1 vccd1 vccd1 final_design.reqhand.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13029_ clknet_leaf_4_clk _00260_ net1098 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08889__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14221__1290 vssd1 vssd1 vccd1 vccd1 _14221__1290/HI net1290 sky130_fd_sc_hd__conb_1
Xfanout1060 final_design.VGA_adr\[10\] vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__buf_2
Xfanout1071 final_design.reqhand.current_client\[3\] vssd1 vssd1 vccd1 vccd1 net1071
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1083 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_4
Xfanout1093 net1094 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08570_ net614 net528 _03517_ net531 vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__o211a_2
XFILLER_0_89_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09370__A _04286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07521_ _01631_ _02471_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07849__C1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11405__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07452_ final_design.cpu.reg_window\[192\] final_design.cpu.reg_window\[224\] net943
+ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06403_ final_design.CPU_instr_adr\[29\] vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07383_ final_design.cpu.reg_window\[258\] final_design.cpu.reg_window\[290\] net947
+ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ net1007 net1003 vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_44_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08813__A1 final_design.CPU_instr_adr\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12070__B1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09053_ net258 _03981_ net1028 vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_96_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout212_A _05951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11140__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ final_design.cpu.reg_window\[720\] final_design.cpu.reg_window\[752\] net879
+ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12782__13 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__inv_2
XFILLER_0_130_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold510 final_design.cpu.reg_window\[814\] vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold521 final_design.cpu.reg_window\[602\] vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 final_design.cpu.reg_window\[695\] vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12373__A1 net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold543 final_design.cpu.reg_window\[235\] vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12670__S net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold554 final_design.cpu.reg_window\[383\] vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap262 _03585_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
Xhold565 final_design.cpu.reg_window\[146\] vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1121_A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold576 final_design.cpu.reg_window\[755\] vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1219_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 final_design.cpu.reg_window\[653\] vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 net160 vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11794__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09955_ _03488_ _04087_ _04873_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout581_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12125__A1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout679_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net633 _03848_ _03849_ _03850_ net259 vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__a311o_1
X_09886_ net265 _04793_ _04803_ _04804_ net451 vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a32o_2
XANTENNA__13540__RESET_B net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1210 final_design.VGA_adr\[1\] vssd1 vssd1 vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 final_design.uart.BAUD_counter\[21\] vssd1 vssd1 vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08837_ final_design.CPU_instr_adr\[10\] final_design.CPU_instr_adr\[9\] _03787_
+ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout846_A net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07552__A1 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08768_ _03713_ _03718_ _03712_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__a21o_1
XANTENNA__12428__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07719_ net610 _02668_ _02643_ net560 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__o211a_1
XANTENNA__11636__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08699_ _02510_ _03647_ _03649_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__nand3_2
XFILLER_0_94_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10730_ _01382_ _05446_ _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_32_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07004__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10661_ net67 _05382_ _05386_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a21o_1
XANTENNA__11034__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11602__X _06157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07939__S net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12400_ _06098_ net354 net341 net1916 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__a22o_1
X_13380_ clknet_leaf_100_clk _00611_ net1187 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[368\]
+ sky130_fd_sc_hd__dfrtp_1
X_10592_ _05315_ _05318_ _05335_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06843__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ net595 _06262_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__nor2_4
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06910__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12262_ net580 _06191_ net511 net373 net1426 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14001_ clknet_leaf_108_clk _01232_ net1215 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[989\]
+ sky130_fd_sc_hd__dfrtp_1
X_11213_ _04772_ _04786_ net660 vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12193_ net1984 net180 net383 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07466__S1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ net230 net2419 net318 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__mux2_1
XANTENNA__12116__A1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11075_ _01388_ _05790_ _05795_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07218__S1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12667__A2 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ net321 _04395_ _04403_ net320 _04944_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10142__A3 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12419__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09190__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11977_ _06179_ net280 net404 net1564 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__a22o_1
XANTENNA__10400__Y _05183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13716_ clknet_leaf_104_clk _00947_ net1202 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[704\]
+ sky130_fd_sc_hd__dfrtp_1
X_10928_ final_design.CPU_instr_adr\[23\] net1054 net814 vssd1 vssd1 vccd1 vccd1 _05657_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13647_ clknet_leaf_93_clk _00878_ net1225 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[635\]
+ sky130_fd_sc_hd__dfrtp_1
X_10859_ net80 _05568_ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__a21o_1
XFILLER_0_160_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13578_ clknet_leaf_1_clk _00809_ net1076 vssd1 vssd1 vccd1 vccd1 final_design.cpu.reg_window\[566\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12529_ _06191_ net349 net328 net1519 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11158__A2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06989__A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07584__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 net310 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_8
Xfanout319 _04117_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_2
XANTENNA__12107__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ _04183_ _04658_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__nand2_1
X_06952_ final_design.cpu.reg_window\[657\] final_design.cpu.reg_window\[689\] net910
+ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__mux2_1
.ends

