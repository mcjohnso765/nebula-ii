module note_div_table (
	note,
	max
);
	reg _sv2v_0;
	input wire [6:0] note;
	output reg [19:0] max;
	always @(*) begin
		if (_sv2v_0)
			;
		case (note)
			7'h00: max = 20'h00000;
			7'h01: max = 20'h954e9;
			7'h02: max = 20'h8ced5;
			7'h03: max = 20'h85047;
			7'h04: max = 20'h7d8d3;
			7'h05: max = 20'h76814;
			7'h06: max = 20'h6fda9;
			7'h07: max = 20'h69937;
			7'h08: max = 20'h63a68;
			7'h09: max = 20'h5e0eb;
			7'h0a: max = 20'h58c74;
			7'h0b: max = 20'h53cbb;
			7'h0c: max = 20'h4f17b;
			7'h0d: max = 20'h4aa75;
			7'h0e: max = 20'h4676a;
			7'h0f: max = 20'h42823;
			7'h10: max = 20'h3ec6a;
			7'h11: max = 20'h3b40a;
			7'h12: max = 20'h37ed5;
			7'h13: max = 20'h34c9b;
			7'h14: max = 20'h31d34;
			7'h15: max = 20'h2f076;
			7'h16: max = 20'h2c63a;
			7'h17: max = 20'h29e5e;
			7'h18: max = 20'h278be;
			7'h19: max = 20'h2553a;
			7'h1a: max = 20'h233b5;
			7'h1b: max = 20'h21412;
			7'h1c: max = 20'h1f635;
			7'h1d: max = 20'h1da05;
			7'h1e: max = 20'h1bf6a;
			7'h1f: max = 20'h1a64e;
			7'h20: max = 20'h18e9a;
			7'h21: max = 20'h1783b;
			7'h22: max = 20'h1631d;
			7'h23: max = 20'h14f2f;
			7'h24: max = 20'h13c5f;
			7'h25: max = 20'h12a9d;
			7'h26: max = 20'h119db;
			7'h27: max = 20'h10a09;
			7'h28: max = 20'h0fb1a;
			7'h29: max = 20'h0ed03;
			7'h2a: max = 20'h0dfb5;
			7'h2b: max = 20'h0d327;
			7'h2c: max = 20'h0c74d;
			7'h2d: max = 20'h0bc1d;
			7'h2e: max = 20'h0b18f;
			7'h2f: max = 20'h0a797;
			7'h30: max = 20'h09e2f;
			7'h31: max = 20'h0954f;
			7'h32: max = 20'h08ced;
			7'h33: max = 20'h08504;
			7'h34: max = 20'h07d8d;
			7'h35: max = 20'h07681;
			7'h36: max = 20'h06fdb;
			7'h37: max = 20'h06993;
			7'h38: max = 20'h063a7;
			7'h39: max = 20'h05e0f;
			7'h3a: max = 20'h058c7;
			7'h3b: max = 20'h053cc;
			7'h3c: max = 20'h04f18;
			7'h3d: max = 20'h04aa7;
			7'h3e: max = 20'h04677;
			7'h3f: max = 20'h04282;
			7'h40: max = 20'h03ec7;
			7'h41: max = 20'h03b41;
			7'h42: max = 20'h037ed;
			7'h43: max = 20'h034ca;
			7'h44: max = 20'h031d3;
			7'h45: max = 20'h02f07;
			7'h46: max = 20'h02c64;
			7'h47: max = 20'h029e6;
			7'h48: max = 20'h0278c;
			7'h49: max = 20'h02554;
			7'h4a: max = 20'h0233b;
			7'h4b: max = 20'h02141;
			7'h4c: max = 20'h01f63;
			7'h4d: max = 20'h01da0;
			7'h4e: max = 20'h01bf7;
			7'h4f: max = 20'h01a65;
			7'h50: max = 20'h018ea;
			7'h51: max = 20'h01784;
			7'h52: max = 20'h01632;
			7'h53: max = 20'h014f3;
			7'h54: max = 20'h013c6;
			7'h55: max = 20'h012aa;
			7'h56: max = 20'h0119e;
			7'h57: max = 20'h010a1;
			7'h58: max = 20'h00fb2;
			7'h59: max = 20'h00ed0;
			7'h5a: max = 20'h00dfb;
			7'h5b: max = 20'h00d32;
			7'h5c: max = 20'h00c75;
			7'h5d: max = 20'h00bc2;
			7'h5e: max = 20'h00b19;
			7'h5f: max = 20'h00a79;
			7'h60: max = 20'h009e3;
			7'h61: max = 20'h00955;
			7'h62: max = 20'h008cf;
			7'h63: max = 20'h00850;
			7'h64: max = 20'h007d9;
			7'h65: max = 20'h00768;
			7'h66: max = 20'h006fe;
			7'h67: max = 20'h00699;
			7'h68: max = 20'h0063a;
			7'h69: max = 20'h005e1;
			7'h6a: max = 20'h0058c;
			7'h6b: max = 20'h0053d;
			7'h6c: max = 20'h004f1;
			7'h6d: max = 20'h004aa;
			7'h6e: max = 20'h00467;
			7'h6f: max = 20'h00428;
			7'h70: max = 20'h003ec;
			7'h71: max = 20'h003b4;
			7'h72: max = 20'h0037f;
			7'h73: max = 20'h0034d;
			7'h74: max = 20'h0031d;
			7'h75: max = 20'h002f0;
			7'h76: max = 20'h002c6;
			7'h77: max = 20'h0029e;
			7'h78: max = 20'h00279;
			7'h79: max = 20'h00255;
			7'h7a: max = 20'h00234;
			7'h7b: max = 20'h00214;
			7'h7c: max = 20'h001f6;
			7'h7d: max = 20'h001da;
			7'h7e: max = 20'h001bf;
			7'h7f: max = 20'h001a6;
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
