* NGSPICE file created from team_06.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

.subckt team_06 clk en gpio_in[0] gpio_in[10] gpio_in[11] gpio_in[12] gpio_in[13]
+ gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17] gpio_in[18] gpio_in[19] gpio_in[1]
+ gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23] gpio_in[24] gpio_in[25] gpio_in[26]
+ gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2] gpio_in[30] gpio_in[31] gpio_in[32]
+ gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3]
+ gpio_oeb[4] gpio_oeb[5] gpio_oeb[6] gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0]
+ gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16]
+ gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22]
+ gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29]
+ gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4]
+ gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XANTENNA__13855__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10669__A1 game.CPU.applesa.ab.absxs.body_x\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_335_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09671_ net1110 _03246_ game.CPU.applesa.ab.absxs.body_y\[36\] net895 _03913_ vssd1
+ vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__a221o_1
XANTENNA__10669__B2 game.CPU.applesa.ab.absxs.body_x\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11119__B net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17202__A2_N net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18869_ clknet_leaf_0_clk _01260_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13174__X _07048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__B game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18895__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10958__B net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_351_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14150__B1_N _07755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16557__B1 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10974__A game.CPU.applesa.ab.absxs.body_x\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1071_A game.CPU.applesa.x\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_335_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09105_ game.CPU.applesa.ab.absxs.body_y\[16\] vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout215_X net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1336_A net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_300_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09036_ game.CPU.applesa.ab.absxs.body_x\[119\] vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19520__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16380__B _02357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout796_A game.CPU.applesa.ab.check_walls.above.walls\[119\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13496__S net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_300_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold340 game.writer.tracker.frame\[243\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_248_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold351 game.writer.tracker.frame\[333\] vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_X net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold362 game.writer.tracker.frame\[89\] vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17285__A1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold373 game.writer.tracker.frame\[265\] vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16088__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold384 game.writer.tracker.frame\[66\] vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_X clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09275__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold395 game.writer.tracker.frame\[92\] vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 game.CPU.applesa.ab.check_walls.above.walls\[47\] vssd1 vssd1 vccd1 vccd1
+ net820 sky130_fd_sc_hd__clkbuf_4
XANTENNA__19670__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout831 game.CPU.applesa.ab.check_walls.above.walls\[7\] vssd1 vssd1 vccd1 vccd1
+ net831 sky130_fd_sc_hd__clkbuf_4
Xfanout842 _06574_ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_4
X_09938_ net1118 net1120 vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__and2_2
XANTENNA__13846__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_183_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout864 net865 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout75_A net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17037__A1 _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout875 net876 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_4
XFILLER_0_245_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15724__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11029__B net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout886 _03368_ vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_125_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09869_ net1085 _03257_ game.CPU.applesa.ab.absxs.body_x\[110\] net923 vssd1 vssd1
+ vccd1 vccd1 _04112_ sky130_fd_sc_hd__a22o_1
Xfanout897 net898 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_4
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_300_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12700__Y _06574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11900_ _05412_ _05785_ _05786_ _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__or4_1
X_12880_ game.writer.tracker.frame\[46\] game.writer.tracker.frame\[47\] net1002 vssd1
+ vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_222_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11831_ _03446_ _05599_ _05607_ _05714_ _05718_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__a311o_1
XANTENNA__11609__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14271__B2 game.CPU.applesa.ab.absxs.body_y\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15740__A game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14550_ _03488_ _04256_ _08419_ vssd1 vssd1 vccd1 vccd1 _08420_ sky130_fd_sc_hd__or3_1
XFILLER_0_261_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ net749 _05265_ _05267_ net570 vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__16555__B _02403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13501_ net224 _07297_ _07374_ net281 vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__o211a_1
X_10713_ _03340_ net425 vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__nor2_1
XANTENNA__19050__CLK net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14481_ _08245_ _08247_ _08249_ _08335_ vssd1 vssd1 vccd1 vccd1 _08355_ sky130_fd_sc_hd__o31a_1
X_11693_ _05567_ _05576_ _05577_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_194_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14023__B2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16220_ _06860_ _02229_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__nor2_2
XFILLER_0_180_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13432_ net693 _06966_ _07305_ net501 vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__o211a_1
XANTENNA__18618__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_354_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_299_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10644_ net1080 _03243_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__nor2_1
XFILLER_0_341_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_311_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16151_ _01741_ _01748_ _02109_ _02162_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_12_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13363_ net502 _07236_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__or2_1
X_10575_ net936 game.CPU.applesa.ab.absxs.body_x\[102\] _04657_ _04660_ vssd1 vssd1
+ vccd1 vccd1 _01153_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15102_ net1203 net1231 game.CPU.applesa.ab.check_walls.above.walls\[130\] vssd1
+ vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__and3_1
X_12314_ _06139_ _06140_ _06150_ _06186_ _06101_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_121_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16082_ net790 net450 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__nor2_1
X_13294_ net231 _07165_ net279 vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__a21o_1
XANTENNA__16720__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16290__B _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18768__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13534__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19910_ clknet_leaf_22_clk game.writer.tracker.next_frame\[505\] net1337 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[505\] sky130_fd_sc_hd__dfrtp_1
X_15033_ net1225 net1256 game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1
+ vccd1 vccd1 _00253_ sky130_fd_sc_hd__and3_1
X_12245_ _05873_ _06130_ _05870_ _05871_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__or4bb_1
XANTENNA__14091__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_clk_X clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17276__A1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_283_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19841_ clknet_leaf_36_clk game.writer.tracker.next_frame\[436\] net1353 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[436\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_254_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12176_ net805 net288 net293 game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1
+ vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_247_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_225_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15474__X net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15915__A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ game.CPU.applesa.ab.absxs.body_x\[16\] net324 vssd1 vssd1 vccd1 vccd1 _05017_
+ sky130_fd_sc_hd__nand2_1
X_16984_ _02465_ net89 _02666_ net2014 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[328\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13298__C1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19772_ clknet_leaf_29_clk game.writer.tracker.next_frame\[367\] net1285 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[367\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_235_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17028__A1 _02369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_322_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11058_ _04943_ _04945_ _04946_ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__or4_1
X_15935_ _03445_ net346 net459 game.CPU.applesa.ab.check_walls.above.walls\[123\]
+ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a22o_1
X_18723_ clknet_leaf_63_clk _01140_ _00460_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[97\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15634__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12610__Y _06487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19390__Q game.CPU.applesa.ab.snake_head_x\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17579__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ _04216_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__inv_2
XANTENNA__16449__C _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18654_ clknet_leaf_51_clk _01071_ _00391_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[68\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15866_ _03322_ net334 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14817_ game.CPU.randy.counter1.count\[13\] game.CPU.randy.counter1.count\[12\] _08619_
+ game.CPU.randy.counter1.count\[14\] vssd1 vssd1 vccd1 vccd1 _08625_ sky130_fd_sc_hd__a31o_1
X_17605_ game.CPU.kyle.L1.cnt_20ms\[6\] _03003_ _03008_ game.CPU.kyle.L1.cnt_20ms\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__a31o_1
X_18585_ clknet_leaf_60_clk _01005_ _00322_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[50\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_235_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15797_ game.CPU.applesa.ab.absxs.body_y\[50\] net441 vssd1 vssd1 vccd1 vccd1 _01809_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__13696__S0 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14262__B2 game.CPU.applesa.ab.absxs.body_x\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_171_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10497__C net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_294_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17536_ _02910_ _02912_ _02918_ _02962_ _04612_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14748_ game.CPU.randy.counter1.count1\[15\] _08571_ vssd1 vssd1 vccd1 vccd1 _08573_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_28_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_318_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_236_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_317_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17467_ _02894_ _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14679_ _08513_ _08514_ _08517_ vssd1 vssd1 vccd1 vccd1 _08518_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_314_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16418_ net235 _02325_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__nor2_1
XFILLER_0_251_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19206_ clknet_leaf_70_clk _00085_ _00854_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.YMAX\[0\]
+ sky130_fd_sc_hd__dfstp_4
XTAP_TAPCELL_ROW_158_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_345_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17398_ game.CPU.kyle.L1.nextState\[3\] game.CPU.kyle.L1.nextState\[2\] _02816_ vssd1
+ vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__or3_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13773__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19137_ net1187 _00179_ _00808_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[182\]
+ sky130_fd_sc_hd__dfrtp_4
X_16349_ _02257_ _02335_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__or2_2
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19068_ net1186 _00103_ _00739_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[113\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15809__B net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_313_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18019_ net660 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__inv_2
XANTENNA__19693__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_247_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout105 net106 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_2
Xfanout116 net118 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__buf_1
XFILLER_0_238_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12233__B net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout127 net128 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_4
Xfanout138 net139 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_2
Xfanout149 net151 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_169_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12801__X _06675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18201__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14486__D1 _08117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_226_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09823__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09723_ net1144 game.CPU.applesa.ab.absxs.body_y\[85\] vssd1 vssd1 vccd1 vccd1 _03966_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__18909__Q game.CPU.applesa.ab.absxs.body_y\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__A game.CPU.applesa.ab.absxs.body_y\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09901__C1 _03981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ net1106 _03469_ _03470_ net1099 vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__a22o_1
XANTENNA__10511__B1 _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_336_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19073__CLK net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09585_ net1103 game.CPU.applesa.ab.check_walls.above.walls\[17\] vssd1 vssd1 vccd1
+ vccd1 _03828_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout165_X net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_43_Left_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout544_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1286_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_355_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_258_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_308_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18644__Q game.CPU.applesa.ab.absxs.body_y\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14005__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14005__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1074_X net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_311_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18910__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09432__A1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16391__A _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14904__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1241_X net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14308__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10360_ game.CPU.walls.rand_wall.counter2\[1\] game.CPU.walls.rand_wall.counter2\[0\]
+ _04519_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_249_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_347_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15719__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Left_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13516__B1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ game.CPU.applesa.ab.absxs.body_x\[67\] vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__inv_2
XANTENNA__11790__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10291_ net1996 _04473_ _04478_ game.CPU.applesa.ab.start_enable vssd1 vssd1 vccd1
+ vccd1 _01315_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_269_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13611__S0 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17258__A1 _02275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12030_ _05912_ _05913_ _05914_ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__or4_1
XFILLER_0_236_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold170 game.writer.tracker.frame\[303\] vssd1 vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09735__A2 game.CPU.applesa.ab.absxs.body_x\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold181 game.writer.tracker.frame\[475\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 game.writer.tracker.frame\[296\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12143__B net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_298_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18111__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_31_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout650 net651 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_4
Xfanout661 net670 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__buf_4
XANTENNA__09733__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_244_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout672 _07401_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15454__B _01454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18819__Q game.CPU.applesa.clk_body vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11982__B net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout683 net692 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_260_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13981_ net952 net828 vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__or2_1
Xfanout694 net695 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__clkbuf_2
XANTENNA__19416__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10879__A game.CPU.applesa.ab.apple_possible\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15720_ game.CPU.applesa.ab.absxs.body_y\[53\] net337 vssd1 vssd1 vccd1 vccd1 _01732_
+ sky130_fd_sc_hd__nand2_1
X_12932_ _06710_ _06712_ net688 vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__mux2_1
XANTENNA__17950__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_358_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_358_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _03468_ net336 vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11046__Y _04936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12863_ game.writer.tracker.frame\[262\] game.writer.tracker.frame\[263\] net996
+ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16566__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14602_ game.CPU.clock1.counter\[5\] _08458_ net268 vssd1 vssd1 vccd1 vccd1 _08459_
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_142_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ net596 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
X_11814_ net825 net312 vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19566__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15582_ game.CPU.applesa.ab.check_walls.above.walls\[91\] net460 net335 _03430_ vssd1
+ vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a2bb2o_1
X_12794_ net493 _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__or2_1
XANTENNA__13452__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17321_ net2021 net732 _02762_ _02422_ _02275_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[569\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__19299__D net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14533_ game.writer.control.current\[1\] game.writer.control.current\[0\] vssd1 vssd1
+ vccd1 vccd1 _08407_ sky130_fd_sc_hd__and2b_1
XFILLER_0_83_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10805__A1 game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11745_ game.CPU.applesa.ab.check_walls.above.walls\[156\] net391 _05630_ _05527_
+ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__o211a_1
XANTENNA__09671__A1 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14086__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09671__B2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11503__A game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17252_ net135 net70 _02280_ net718 vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__o31a_1
X_14464_ game.CPU.applesa.ab.absxs.body_x\[60\] net1075 vssd1 vssd1 vccd1 vccd1 _08338_
+ sky130_fd_sc_hd__xor2_1
X_11676_ game.CPU.applesa.ab.check_walls.above.walls\[127\] net258 _05560_ _05564_
+ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__o211a_2
XFILLER_0_153_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13755__A0 game.writer.tracker.frame\[161\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16203_ _01684_ _01685_ _01687_ _01688_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a22o_1
X_13415_ net240 _07271_ _07288_ _06860_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_221_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18590__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11222__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17183_ _02487_ net74 _02726_ net1694 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[467\]
+ sky130_fd_sc_hd__a22o_1
X_10627_ game.CPU.applesa.ab.absxs.body_x\[59\] net327 _04681_ net933 vssd1 vssd1
+ vccd1 vccd1 _01122_ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14395_ game.CPU.applesa.ab.absxs.body_y\[71\] net946 vssd1 vssd1 vccd1 vccd1 _08269_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_3_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16134_ game.CPU.applesa.ab.absxs.body_y\[22\] net440 net469 game.CPU.applesa.ab.absxs.body_x\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a2bb2o_1
X_13346_ net702 _06617_ _07219_ net226 vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_231_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09908__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10558_ game.CPU.applesa.ab.absxs.body_x\[23\] _04645_ _04652_ game.CPU.applesa.ab.absxs.body_x\[19\]
+ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11781__A2 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16065_ game.CPU.applesa.ab.check_walls.above.walls\[196\] net450 vssd1 vssd1 vccd1
+ vccd1 _02077_ sky130_fd_sc_hd__xnor2_1
X_13277_ net694 _07150_ _07147_ net220 vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__o211a_1
XANTENNA__13602__S0 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489_ net1117 _04578_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__or2_2
XANTENNA__17249__A1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15016_ net1220 net1248 game.CPU.applesa.ab.check_walls.above.walls\[44\] vssd1 vssd1
+ vccd1 vccd1 _00235_ sky130_fd_sc_hd__and3_1
X_12228_ net809 net417 _05961_ _05962_ _06113_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11533__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19824_ clknet_leaf_39_clk game.writer.tracker.next_frame\[419\] net1352 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[419\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15645__A game.CPU.applesa.ab.check_walls.above.walls\[74\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12159_ _06043_ _06044_ _06045_ _06042_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__a211o_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19755_ clknet_leaf_25_clk game.writer.tracker.next_frame\[350\] net1321 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[350\] sky130_fd_sc_hd__dfrtp_1
X_16967_ _02429_ net96 _02660_ net1742 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[317\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_316_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_263_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_264_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18706_ clknet_leaf_50_clk _01123_ _00443_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[64\]
+ sky130_fd_sc_hd__dfrtp_4
X_15918_ net793 net342 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__nand2_1
XANTENNA__12494__B1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19686_ clknet_leaf_34_clk game.writer.tracker.next_frame\[281\] net1319 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[281\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_242_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16898_ _02300_ net92 _02641_ net1853 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[267\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19909__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16224__A2 net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18637_ clknet_leaf_61_clk _01054_ _00374_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_15849_ game.CPU.applesa.ab.absxs.body_y\[99\] net432 vssd1 vssd1 vccd1 vccd1 _01861_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__16476__A _02289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09370_ net916 game.CPU.applesa.ab.check_walls.above.walls\[33\] game.CPU.applesa.ab.check_walls.above.walls\[35\]
+ net926 _03612_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__a221o_1
XANTENNA__13443__C1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18568_ clknet_leaf_8_clk _00988_ _00305_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17519_ _02844_ _02924_ _02946_ _02921_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a211o_1
XFILLER_0_191_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18499_ net586 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__inv_2
XANTENNA__18933__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09662__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12509__A game.CPU.applesa.ab.absxs.body_x\[73\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12892__S1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09662__B2 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_306_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_305_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16482__Y _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload64_A clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11132__B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout125_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10971__B net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14443__B net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10575__A3 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12244__A game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1034_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout494_A _06596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19439__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1201_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10732__B1 _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_342_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09706_ net1094 _03412_ _03944_ _03946_ _03948_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a2111o_1
XANTENNA__19589__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19537__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11307__B net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09637_ _03872_ _03873_ _03874_ _03879_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__or4_2
XFILLER_0_179_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16386__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout547_X net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09568_ net904 game.CPU.applesa.ab.absxs.body_y\[78\] _03302_ net1158 vssd1 vssd1
+ vccd1 vccd1 _03811_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09837__A1_N net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_104_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17176__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09499_ net1139 net819 vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11530_ net821 net257 vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_322_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16923__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11042__B net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11461_ game.CPU.applesa.ab.check_walls.above.walls\[18\] net768 vssd1 vssd1 vccd1
+ vccd1 _05350_ sky130_fd_sc_hd__xor2_2
XFILLER_0_80_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_311_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13200_ game.writer.tracker.frame\[396\] game.writer.tracker.frame\[397\] net1020
+ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__mux2_1
Xwire358 _07875_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_1
XFILLER_0_296_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10412_ game.CPU.randy.f1.state\[1\] _03222_ _04558_ vssd1 vssd1 vccd1 vccd1 _04559_
+ sky130_fd_sc_hd__a21oi_1
X_11392_ net805 net257 vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__or2_1
XANTENNA__09728__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14180_ game.CPU.applesa.ab.absxs.body_x\[17\] net1063 vssd1 vssd1 vccd1 vccd1 _08054_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13131_ _07001_ _07003_ net679 vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__mux2_1
X_10343_ net1809 _04505_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__nor2_1
XANTENNA__17945__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13062_ game.writer.tracker.frame\[242\] game.writer.tracker.frame\[243\] net1027
+ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__mux2_1
X_10274_ net1170 _04362_ _04375_ net1172 vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__o22a_1
XFILLER_0_249_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_280_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11515__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net811 net298 net291 net812 vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__a22o_1
XANTENNA__11993__A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17870_ _03185_ _03188_ _03189_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_306_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09463__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16821_ _02513_ net100 _02606_ net2027 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[225\]
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__19960__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_144_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout480 net486 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__buf_2
XANTENNA__15662__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout491 net493 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_4
X_19540_ clknet_leaf_33_clk game.writer.tracker.next_frame\[135\] net1296 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[135\] sky130_fd_sc_hd__dfrtp_1
X_16752_ net164 _02396_ net110 _02585_ game.writer.tracker.frame\[176\] vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.next_frame\[176\] sky130_fd_sc_hd__a32o_1
XFILLER_0_283_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13964_ net882 game.CPU.applesa.ab.check_walls.above.walls\[177\] game.CPU.applesa.ab.check_walls.above.walls\[182\]
+ net855 vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_205_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09877__D1 _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15703_ _03462_ net332 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__xnor2_1
X_12915_ _06674_ _06677_ net683 vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19471_ clknet_leaf_19_clk game.writer.tracker.next_frame\[66\] net1335 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[66\] sky130_fd_sc_hd__dfrtp_1
X_16683_ _02252_ _02257_ net98 net718 vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__o31a_1
XANTENNA__15912__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11217__B net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18956__CLK net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13895_ net878 game.CPU.applesa.ab.check_walls.above.walls\[58\] _03413_ net985 vssd1
+ vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_204_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15634_ game.CPU.applesa.ab.absxs.body_y\[83\] net431 vssd1 vssd1 vccd1 vccd1 _01646_
+ sky130_fd_sc_hd__xnor2_1
X_18422_ net626 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
X_12846_ game.writer.tracker.frame\[312\] game.writer.tracker.frame\[313\] net1033
+ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_291_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ net593 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__inv_2
X_15565_ _03363_ _06545_ _06548_ _01583_ vssd1 vssd1 vccd1 vccd1 game.writer.updater.update.next\[0\]
+ sky130_fd_sc_hd__a31o_1
X_12777_ game.writer.tracker.frame\[126\] game.writer.tracker.frame\[127\] net1033
+ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__mux2_1
XANTENNA__09644__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16509__A3 _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09644__B2 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17304_ game.writer.tracker.frame\[557\] net722 _02757_ vssd1 vssd1 vccd1 vccd1 _02758_
+ sky130_fd_sc_hd__and3_1
XANTENNA__11233__A game.CPU.applesa.ab.absxs.body_x\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14516_ _08382_ _08383_ _08385_ _08387_ vssd1 vssd1 vccd1 vccd1 _08390_ sky130_fd_sc_hd__or4_1
X_11728_ _05610_ _05614_ _05615_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__and3_1
X_18284_ net621 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
XFILLER_0_232_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15496_ net883 _01505_ _01507_ net865 _01519_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17235_ net154 _02423_ net79 _02739_ net1595 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[506\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14447_ game.CPU.applesa.ab.absxs.body_x\[89\] net882 net947 _03326_ vssd1 vssd1
+ vccd1 vccd1 _08321_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ net830 net317 vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__nand2_1
XFILLER_0_303_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18016__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17166_ _02460_ net122 net121 _02722_ net1559 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[454\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11887__B net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14378_ _03330_ net958 net938 _03328_ vssd1 vssd1 vccd1 vccd1 _08252_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12335__Y game.CPU.applesa.twoapples.absxs.next_head\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16117_ _03303_ net334 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11754__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13329_ net219 _07200_ _07202_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__a21o_1
X_17097_ game.writer.tracker.frame\[407\] _02700_ vssd1 vssd1 vccd1 vccd1 _02701_
+ sky130_fd_sc_hd__and2_1
XANTENNA__16142__A1 game.CPU.applesa.ab.absxs.body_y\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15078__C game.CPU.applesa.ab.check_walls.above.walls\[106\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16142__B2 game.CPU.applesa.ab.absxs.body_y\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_3_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_16048_ _02052_ _02055_ _02058_ _02059_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_94_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12703__A1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13447__X _07321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_244_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19807_ clknet_leaf_37_clk game.writer.tracker.next_frame\[402\] net1354 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[402\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19731__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17999_ net637 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__inv_2
XFILLER_0_208_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19738_ clknet_leaf_18_clk game.writer.tracker.next_frame\[333\] net1289 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[333\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16477__Y _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09660__X _03903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_239_Right_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11127__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19669_ clknet_leaf_30_clk game.writer.tracker.next_frame\[264\] net1292 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[264\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09883__A1 _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19881__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09422_ _03658_ _03659_ _03660_ _03661_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__or4_1
XFILLER_0_126_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14438__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09353_ net1102 _03291_ game.CPU.applesa.ab.absxs.body_y\[8\] net893 vssd1 vssd1
+ vccd1 vccd1 _03596_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_255_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout242_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12239__A game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12865__S1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11143__A game.CPU.applesa.ab.absxs.body_y\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_129_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11442__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09284_ net756 _03527_ net755 net1732 vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11165__A2_N net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1151_A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout128_X net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1249_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09548__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14392__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14173__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19261__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11745__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_344_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16133__B2 game.CPU.applesa.ab.absxs.body_y\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1037_X net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18829__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12096__A1_N net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_266_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10705__B1 _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09571__B1 game.CPU.applesa.ab.absxs.body_y\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18979__CLK net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ game.CPU.applesa.ab.absxs.body_x\[29\] vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__inv_2
XFILLER_0_215_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16987__A3 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11318__A _05194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16828__B net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15732__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10961_ game.CPU.applesa.ab.absxs.body_y\[119\] net398 vssd1 vssd1 vccd1 vccd1 _04851_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_355_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_206_Right_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14188__X _08062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net1004 net969 vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__nand2_4
XANTENNA__16547__C _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ net476 _07551_ _07552_ _07553_ net201 vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__a311o_1
XFILLER_0_195_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10892_ net769 net765 net759 net773 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__or4b_1
XFILLER_0_329_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_277_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10876__B game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14348__B net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12631_ game.CPU.applesa.ab.absxs.body_y\[10\] net519 _03356_ game.CPU.applesa.twoapples.absxs.next_head\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_333_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_219_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12149__A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15350_ game.writer.updater.commands.count\[15\] game.writer.updater.commands.count\[14\]
+ game.writer.updater.commands.count\[13\] vssd1 vssd1 vccd1 vccd1 _08892_ sky130_fd_sc_hd__or3_1
XFILLER_0_182_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12562_ game.CPU.applesa.ab.absxs.body_y\[119\] net366 vssd1 vssd1 vccd1 vccd1 _06439_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ game.CPU.applesa.ab.absxs.body_y\[30\] net949 vssd1 vssd1 vccd1 vccd1 _08175_
+ sky130_fd_sc_hd__xor2_1
X_11513_ game.CPU.applesa.ab.check_walls.above.walls\[0\] net777 vssd1 vssd1 vccd1
+ vccd1 _05402_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19604__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15281_ _08831_ _08834_ vssd1 vssd1 vccd1 vccd1 _08835_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10892__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12493_ game.CPU.applesa.ab.absxs.body_x\[81\] net375 game.CPU.applesa.twoapples.absxs.next_head\[7\]
+ _03328_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__a22o_1
X_17020_ _02579_ _02670_ net717 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__o21a_1
XANTENNA__14383__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14232_ _08100_ _08101_ _08105_ _08097_ vssd1 vssd1 vccd1 vccd1 _08106_ sky130_fd_sc_hd__a211o_1
XFILLER_0_269_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11444_ game.CPU.applesa.ab.check_walls.above.walls\[72\] net779 vssd1 vssd1 vccd1
+ vccd1 _05333_ sky130_fd_sc_hd__xor2_1
XFILLER_0_202_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12933__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ net923 net1057 net965 net899 _08036_ vssd1 vssd1 vccd1 vccd1 _08037_ sky130_fd_sc_hd__a221o_1
XANTENNA__17321__B1 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11375_ _05252_ _05250_ _05251_ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_308_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13114_ net504 _06985_ _06987_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__a21o_1
XANTENNA__19754__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10326_ _04500_ _04503_ vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_150_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15907__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14094_ net1049 game.CPU.applesa.ab.check_walls.above.walls\[11\] vssd1 vssd1 vccd1
+ vccd1 _07968_ sky130_fd_sc_hd__xor2_1
X_18971_ net1199 _00165_ _00642_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__17394__B _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13489__A2 _07144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13045_ net275 _06918_ _06915_ net243 vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__o211a_1
X_17922_ net605 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__inv_2
X_10257_ net779 net771 vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__nor2_2
Xfanout1220 net1221 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__buf_2
XANTENNA__16427__A2 _02310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12161__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1231 net1232 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__dlymetal6s2s_1
X_17853_ game.writer.updater.commands.count\[11\] _03172_ vssd1 vssd1 vccd1 vccd1
+ _03177_ sky130_fd_sc_hd__or2_1
X_10188_ net1168 net773 vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__nand2_1
Xfanout1242 net1257 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_245_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1253 net1254 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_206_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1264 game.CPU.clock1.game_state\[1\] vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__buf_2
X_16804_ _02328_ net144 net99 net728 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__o31a_1
Xfanout1275 game.CPU.speed1.Qa\[1\] vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__buf_2
Xfanout1286 net1293 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__clkbuf_2
Xfanout1297 net1307 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__clkbuf_2
X_17784_ _03126_ game.CPU.applesa.twoapples.count\[3\] game.CPU.applesa.twoapples.count\[1\]
+ game.CPU.applesa.twoapples.count\[2\] vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__and4b_1
X_14996_ net1224 net1255 game.CPU.applesa.ab.check_walls.above.walls\[24\] vssd1 vssd1
+ vccd1 vccd1 _00213_ sky130_fd_sc_hd__and3_1
XANTENNA__16297__Y _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19523_ clknet_leaf_21_clk game.writer.tracker.next_frame\[118\] net1335 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[118\] sky130_fd_sc_hd__dfrtp_1
X_16735_ _02365_ _02561_ net719 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__o21a_1
X_13947_ _07817_ _07818_ _07819_ _07820_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__or4_4
XANTENNA__15642__B net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_319_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16666_ net152 _02431_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__and2_1
X_19454_ clknet_leaf_43_clk game.writer.tracker.next_frame\[49\] net1327 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[49\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09640__B net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19134__CLK net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ net984 _03438_ _03439_ net950 _07751_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__o221a_1
XFILLER_0_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14258__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18405_ net602 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
X_15617_ game.CPU.applesa.ab.check_walls.above.walls\[86\] net333 vssd1 vssd1 vccd1
+ vccd1 _01629_ sky130_fd_sc_hd__or2_1
X_12829_ net162 net173 vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__nand2_1
X_16597_ game.writer.tracker.frame\[97\] _02510_ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__nand2_1
X_19385_ clknet_leaf_3_clk _01391_ _00965_ vssd1 vssd1 vccd1 vccd1 game.CPU.bodymain1.main.score\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_243_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15548_ _01552_ _01568_ _01567_ _01564_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__o211a_1
X_18336_ net599 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14545__Y game.CPU.walls.rand_wall.abduyd.next_wall\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19284__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18742__Q game.CPU.applesa.ab.absxs.body_x\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18267_ net649 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XFILLER_0_343_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15479_ _01502_ _01503_ _01492_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_330_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17218_ _02389_ net142 net119 _02735_ net1592 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[493\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__09368__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18198_ net580 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15089__B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_303_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_250_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12506__B net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17149_ _02424_ net58 _02716_ net1623 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[443\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14126__B1 game.CPU.applesa.ab.check_walls.above.walls\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap455 net456 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_338_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09971_ net1078 _04198_ _04199_ _04156_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__o31a_1
XANTENNA__15817__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_308_Right_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15874__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19811__RESET_B net1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_283_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_354_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16134__A2_N net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13101__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout457_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16367__C _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1199_A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14168__B net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ net1138 game.CPU.applesa.ab.check_walls.above.walls\[134\] vssd1 vssd1 vccd1
+ vccd1 _03648_ sky130_fd_sc_hd__xor2_1
XANTENNA__19627__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout245_X net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout624_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_338_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09336_ net1090 game.CPU.applesa.ab.absxs.body_x\[90\] vssd1 vssd1 vccd1 vccd1 _03579_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12612__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_350_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ game.CPU.randy.counter1.count1\[2\] vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12256__X _06142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14184__A game.CPU.applesa.ab.absxs.body_y\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1154_X net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11601__A game.CPU.applesa.ab.check_walls.above.walls\[98\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18651__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19777__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ game.CPU.applesa.ab.check_walls.above.walls\[128\] vssd1 vssd1 vccd1 vccd1
+ _03447_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout993_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12416__B game.CPU.applesa.twoapples.absxs.next_head\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_214_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14471__X _08345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16657__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16830__C net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14117__B1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ game.CPU.applesa.ab.absxs.body_y\[51\] net397 vssd1 vssd1 vccd1 vccd1 _05050_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_248_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15727__B net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_286_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout879_X net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ _04315_ net1463 _04311_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__mux2_1
X_11091_ game.CPU.applesa.ab.absxs.body_x\[58\] net409 vssd1 vssd1 vccd1 vccd1 _04981_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10651__S _04690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13340__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10042_ net1174 _04226_ _04237_ net1170 vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__o22a_1
XANTENNA__12774__S0 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16398__X _02370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold30 game.CPU.reset_button1.eD1.Q2 vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12151__B net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold41 game.CPU.applesa.twomode.number\[0\] vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_303_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17082__A2 _02693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold52 game.CPU.kyle.L1.lcd_rs vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ game.CPU.randy.f1.c1.count\[9\] _08643_ vssd1 vssd1 vccd1 vccd1 _08645_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout60_X net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold63 game.CPU.applesa.apple_location2_n\[1\] vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19157__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold74 net41 vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 game.writer.tracker.frame\[458\] vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13801_ game.writer.tracker.frame\[423\] net711 net674 game.writer.tracker.frame\[424\]
+ vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__o22a_1
Xhold96 game.writer.tracker.frame\[45\] vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09741__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_349_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14781_ _03516_ net139 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__and2_1
XFILLER_0_242_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11993_ net826 net553 vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__or2_1
XANTENNA__13643__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14359__A game.CPU.applesa.ab.absxs.body_y\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16520_ net190 net125 _02460_ _02459_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[70\]
+ sky130_fd_sc_hd__a31o_1
X_13732_ game.writer.tracker.frame\[219\] net710 net673 game.writer.tracker.frame\[220\]
+ vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__o22a_1
XFILLER_0_202_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10944_ game.CPU.applesa.ab.absxs.body_x\[28\] net416 vssd1 vssd1 vccd1 vccd1 _04834_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_329_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16451_ net206 _02326_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__nor2_8
XFILLER_0_85_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13663_ _07535_ _07536_ net483 vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__mux2_1
X_10875_ _04775_ _04776_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16593__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16574__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_329_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15402_ game.writer.updater.commands.count\[15\] _01429_ game.writer.updater.commands.count\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_197_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19170_ clknet_leaf_58_clk _00288_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.collisions
+ sky130_fd_sc_hd__dfxtp_1
X_12614_ _06489_ _06456_ _06488_ _06490_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__and4b_2
X_16382_ _02274_ _02359_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__or2_1
XANTENNA__11610__A2_N net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ game.writer.tracker.frame\[381\] game.writer.tracker.frame\[383\] game.writer.tracker.frame\[384\]
+ game.writer.tracker.frame\[382\] net979 net1032 vssd1 vssd1 vccd1 vccd1 _07468_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13800__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18121_ net577 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__inv_2
XFILLER_0_344_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_314_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15333_ game.CPU.applesa.twomode.number\[3\] _08871_ vssd1 vssd1 vccd1 vccd1 _08876_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__11957__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18562__Q game.CPU.applesa.ab.absxs.body_y\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12545_ game.CPU.applesa.ab.absxs.body_x\[40\] net384 _06420_ _06421_ vssd1 vssd1
+ vccd1 vccd1 _06422_ sky130_fd_sc_hd__o211a_1
XFILLER_0_325_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14094__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18052_ net656 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11511__A game.CPU.applesa.ab.check_walls.above.walls\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15264_ _01263_ _08818_ vssd1 vssd1 vccd1 vccd1 _08820_ sky130_fd_sc_hd__nor2_1
XFILLER_0_352_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12476_ game.CPU.applesa.ab.absxs.body_y\[31\] net364 vssd1 vssd1 vccd1 vccd1 _06353_
+ sky130_fd_sc_hd__xnor2_1
X_17003_ _02489_ net83 _02672_ net1903 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[341\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11230__B net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ game.CPU.applesa.ab.absxs.body_x\[93\] net881 net959 _03297_ vssd1 vssd1
+ vccd1 vccd1 _08089_ sky130_fd_sc_hd__a22o_1
XANTENNA__15918__A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_5 _02179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ net826 net252 vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__or2_1
X_15195_ game.CPU.applesa.normal1.counter_flip game.CPU.applesa.normal1.number\[4\]
+ vssd1 vssd1 vccd1 vccd1 _08765_ sky130_fd_sc_hd__and2b_1
XFILLER_0_300_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16648__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09916__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ _07956_ _07962_ _08017_ _08019_ vssd1 vssd1 vccd1 vccd1 _08020_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_286_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15637__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11358_ game.CPU.applesa.ab.check_walls.above.walls\[140\] net249 vssd1 vssd1 vccd1
+ vccd1 _05247_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10393__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14541__B _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15856__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ _04491_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__inv_2
X_18954_ clknet_leaf_68_clk net1419 _00625_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14077_ net1171 net862 game.CPU.applesa.ab.YMAX\[2\] net852 _07950_ vssd1 vssd1 vccd1
+ vccd1 _07951_ sky130_fd_sc_hd__a221o_1
XANTENNA__09635__B game.CPU.applesa.ab.absxs.body_y\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11289_ _04993_ _05135_ _05137_ _05136_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_33_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13331__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13028_ _06900_ _06901_ net506 vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_265_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17905_ net661 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__inv_2
XFILLER_0_206_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12061__B net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18885_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[15\] _00580_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[15\] sky130_fd_sc_hd__dfrtp_1
Xfanout1050 net1051 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17073__A2 net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13725__X _07599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15653__A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1061 net1062 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_163_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17836_ _03150_ _03163_ _03164_ net182 game.writer.updater.commands.count\[6\] vssd1
+ vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__a32o_1
XFILLER_0_177_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10696__A2 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1072 net1077 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__buf_4
Xfanout1083 net1088 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__buf_6
XANTENNA__16281__B1 _08028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1094 net1095 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__buf_4
XANTENNA__09651__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16820__A2 _02359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09838__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17767_ game.CPU.applesa.twoapples.count_luck\[5\] game.CPU.applesa.twoapples.count_luck\[4\]
+ _03116_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__and3_1
XFILLER_0_324_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09838__B2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ net1226 net1253 game.CPU.applesa.ab.check_walls.above.walls\[7\] vssd1 vssd1
+ vccd1 vccd1 _00154_ sky130_fd_sc_hd__and3_1
XFILLER_0_344_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13190__S0 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19506_ clknet_leaf_29_clk game.writer.tracker.next_frame\[101\] net1283 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[101\] sky130_fd_sc_hd__dfrtp_1
X_16718_ net160 _02289_ _02297_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__and3_2
XFILLER_0_221_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_297_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17698_ game.CPU.walls.rand_wall.count\[0\] net1175 vssd1 vssd1 vccd1 vccd1 _03077_
+ sky130_fd_sc_hd__or2_1
X_19437_ clknet_leaf_39_clk game.writer.tracker.next_frame\[32\] net1332 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[32\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_239_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16649_ net114 net158 _02413_ net730 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16484__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_252_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18674__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19368_ clknet_leaf_71_clk _01374_ _00949_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_09121_ game.CPU.applesa.ab.XMAX\[1\] vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__inv_2
XFILLER_0_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18319_ net615 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_99_Left_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19299_ clknet_leaf_69_clk net408 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.x_final\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12517__A game.CPU.applesa.ab.absxs.body_y\[69\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_127_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11421__A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_343_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09052_ game.CPU.applesa.ab.absxs.body_y\[77\] vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__inv_2
XFILLER_0_303_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold500 game.writer.tracker.frame\[509\] vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12951__S net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10908__A0 net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold511 game.writer.tracker.frame\[327\] vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12804__X _06678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold522 game.writer.tracker.frame\[34\] vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold533 game.CPU.randy.f1.c1.count\[17\] vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16639__A2 _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12373__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__A net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09774__B1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold544 game.writer.tracker.frame\[559\] vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 game.writer.tracker.frame\[352\] vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 game.writer.tracker.frame\[136\] vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14451__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold577 game.writer.tracker.frame\[137\] vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 game.CPU.kyle.L1.cnt_20ms\[10\] vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09545__B game.CPU.applesa.ab.absxs.body_x\[114\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09954_ _03527_ _04158_ game.CPU.bodymain1.main.score\[0\] vssd1 vssd1 vccd1 vccd1
+ _04185_ sky130_fd_sc_hd__a21oi_1
Xhold599 game.writer.tracker.frame\[27\] vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_263_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13322__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_271_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09885_ _04121_ _04122_ _04123_ _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout574_A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout195_X net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17064__A2 _02455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_291_Right_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_271_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16378__B _02289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09561__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16811__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_339_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09829__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09829__B2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11636__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_352_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1271_X net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_274_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10660_ game.CPU.applesa.ab.absxs.body_x\[27\] _04695_ _04698_ game.CPU.applesa.ab.absxs.body_x\[23\]
+ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17119__A3 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13484__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09319_ net900 game.CPU.applesa.ab.absxs.body_y\[65\] game.CPU.applesa.ab.absxs.body_y\[64\]
+ net894 _03558_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__a221o_1
X_10591_ game.CPU.applesa.ab.absxs.body_x\[108\] _04665_ _04666_ game.CPU.applesa.ab.absxs.body_x\[104\]
+ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12427__A game.CPU.applesa.ab.absxs.body_y\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12330_ net1162 _04224_ _06211_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a21o_1
XANTENNA__14338__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16878__A2 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10611__A2 _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11050__B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ game.CPU.applesa.ab.check_walls.above.walls\[166\] net417 vssd1 vssd1 vccd1
+ vccd1 _06147_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12861__S net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_188_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14000_ net877 game.CPU.applesa.ab.check_walls.above.walls\[74\] game.CPU.applesa.ab.check_walls.above.walls\[78\]
+ net855 _07869_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__o221a_1
XANTENNA__12364__A2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ game.CPU.applesa.ab.absxs.body_y\[95\] net396 vssd1 vssd1 vccd1 vccd1 _05102_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__15457__B _01454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12192_ _06074_ _06075_ _06076_ _06077_ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__or4_1
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
Xoutput42 net42 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_339_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11143_ game.CPU.applesa.ab.absxs.body_y\[96\] net537 vssd1 vssd1 vccd1 vccd1 _05033_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13313__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14510__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17672__B _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10127__A1 net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15951_ _01951_ _01952_ _01957_ _01962_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__or4_1
X_11074_ game.CPU.applesa.ab.absxs.body_x\[42\] net410 vssd1 vssd1 vccd1 vccd1 _04964_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__16569__A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10025_ net1090 _04232_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__nand2_1
X_14902_ net1144 _08426_ vssd1 vssd1 vccd1 vccd1 _08679_ sky130_fd_sc_hd__nand2_1
X_15882_ game.CPU.applesa.ab.check_walls.above.walls\[138\] net465 vssd1 vssd1 vccd1
+ vccd1 _01894_ sky130_fd_sc_hd__nor2_1
X_18670_ clknet_leaf_10_clk _01087_ _00407_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[100\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16288__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09471__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16802__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17621_ _03028_ _03029_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__nor2_1
X_14833_ _04332_ _08633_ _08634_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[2\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__13616__A2 game.writer.tracker.frame\[320\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14089__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11506__A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17552_ _08443_ _02782_ net426 vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__and3b_1
XANTENNA__18697__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14764_ game.CPU.randy.counter1.count\[11\] _04356_ _08492_ vssd1 vssd1 vccd1 vccd1
+ _08585_ sky130_fd_sc_hd__and3_1
X_11976_ game.CPU.applesa.ab.apple_possible\[5\] _04775_ vssd1 vssd1 vccd1 vccd1 _05863_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__11627__B2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_316_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19942__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_230_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13715_ net220 _07588_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__or2_1
X_16503_ net219 _02447_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__nor2_2
XANTENNA__11225__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10927_ _03289_ net406 vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15920__B net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17483_ _02883_ _02911_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__nor2_1
XFILLER_0_357_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14695_ game.CPU.randy.counter1.count1\[11\] _08491_ _08525_ _08533_ vssd1 vssd1
+ vccd1 vccd1 _08534_ sky130_fd_sc_hd__a211o_1
X_19222_ clknet_leaf_69_clk _01316_ _00861_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_location\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13646_ game.writer.tracker.frame\[26\] net844 net711 game.writer.tracker.frame\[27\]
+ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__o22a_1
X_16434_ net116 net165 _02396_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10858_ _04739_ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_344_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_317_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16365_ net236 _02264_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_15_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19153_ net1187 _00196_ _00824_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[198\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_143_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13577_ _07449_ _07450_ net511 vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__mux2_1
XANTENNA__12337__A net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10789_ _03341_ net561 vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__nor2_1
X_15316_ game.CPU.applesa.twomode.number\[0\] _08856_ net757 vssd1 vssd1 vccd1 vccd1
+ _08862_ sky130_fd_sc_hd__a21oi_1
X_18104_ net628 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__inv_2
XANTENNA__16869__A2 _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10602__A2 _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12528_ game.CPU.applesa.ab.absxs.body_y\[99\] net364 net529 game.CPU.applesa.ab.absxs.body_x\[99\]
+ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_325_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16296_ _02245_ _02295_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__nand2_1
X_19084_ net1177 _00120_ _00755_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[129\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12480__A1_N game.CPU.applesa.ab.absxs.body_y\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_240_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15247_ _08804_ _08805_ _08806_ _08807_ vssd1 vssd1 vccd1 vccd1 _08808_ sky130_fd_sc_hd__and4_4
X_18035_ net590 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09917__Y _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12459_ _06326_ _06327_ _06329_ _06335_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__or4_2
XFILLER_0_313_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15541__A2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_327_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19322__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13869__A1_N game.CPU.applesa.ab.XMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15178_ _08751_ _08753_ vssd1 vssd1 vccd1 vccd1 _08754_ sky130_fd_sc_hd__nand2_1
XANTENNA__11895__B net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19403__RESET_B net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10366__A1 game.CPU.applesa.ab.absxs.body_y\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11563__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14129_ _07997_ _08001_ _08002_ vssd1 vssd1 vccd1 vccd1 _08003_ sky130_fd_sc_hd__and3_1
XFILLER_0_249_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19986_ clknet_leaf_45_clk _01410_ net1304 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout309 _05606_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__buf_4
XFILLER_0_281_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18937_ clknet_leaf_15_clk net1391 net1282 vssd1 vssd1 vccd1 vccd1 game.CPU.reset_button1.eD1.D
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10118__A1 game.CPU.applesa.enable_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16479__A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10304__B net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19472__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17046__A2 _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09670_ net926 game.CPU.applesa.ab.absxs.body_x\[39\] game.CPU.applesa.ab.absxs.body_x\[36\]
+ net912 vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__a22o_1
XANTENNA__11866__A1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10669__A2 _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18868_ clknet_leaf_0_clk _01259_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17819_ net182 _03151_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__nor2_1
X_18799_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[2\] _00536_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_221_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11416__A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14280__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11135__B net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15830__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16557__B2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout155_A _02270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_335_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10974__B net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_351_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout322_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12247__A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1064_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09104_ game.CPU.applesa.ab.absxs.body_y\[17\] vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__inv_2
XANTENNA__12594__A2 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_304_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15517__C1 _08028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09035_ game.CPU.applesa.ab.absxs.body_x\[16\] vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout110_X net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_300_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1231_A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout208_X net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1329_A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold330 game.writer.tracker.frame\[157\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold341 game.writer.tracker.frame\[173\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold352 game.writer.tracker.frame\[306\] vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 game.writer.tracker.frame\[251\] vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A game.CPU.applesa.ab.check_walls.above.walls\[151\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19815__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold374 game.writer.tracker.frame\[91\] vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17285__A2 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold385 game.writer.tracker.frame\[135\] vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_6_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold396 game.writer.tracker.frame\[511\] vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 game.CPU.applesa.ab.check_walls.above.walls\[84\] vssd1 vssd1 vccd1 vccd1
+ net810 sky130_fd_sc_hd__clkbuf_4
Xfanout821 game.CPU.applesa.ab.check_walls.above.walls\[46\] vssd1 vssd1 vccd1 vccd1
+ net821 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_309_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout832 game.CPU.applesa.ab.check_walls.above.walls\[4\] vssd1 vssd1 vccd1 vccd1
+ net832 sky130_fd_sc_hd__clkbuf_4
X_09937_ net1121 _04172_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__nand2_1
Xfanout843 _06574_ vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__buf_4
XANTENNA_fanout956_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_183_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13365__X _07239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout865 net866 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_6
Xfanout876 _03373_ vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__buf_8
XANTENNA__11857__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09868_ net1149 game.CPU.applesa.ab.absxs.body_y\[109\] vssd1 vssd1 vccd1 vccd1 _04111_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_125_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout887 _03368_ vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__buf_4
Xfanout898 net901 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_6
XANTENNA__11857__B2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_300_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19965__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout68_A _02373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11012__A1_N game.CPU.applesa.ab.absxs.body_x\[53\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09291__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09799_ _04038_ _04040_ _04041_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__nand3b_2
XTAP_TAPCELL_ROW_222_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11326__A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11830_ net571 _05551_ _05552_ net747 _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__a221o_1
XANTENNA__14271__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11045__B net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15740__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout911_X net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ game.CPU.applesa.ab.check_walls.above.walls\[181\] net307 vssd1 vssd1 vccd1
+ vccd1 _05649_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16548__B2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13500_ net482 _07294_ _07296_ net204 vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10712_ game.CPU.applesa.ab.absxs.body_y\[61\] net425 _04712_ net933 vssd1 vssd1
+ vccd1 vccd1 _01068_ sky130_fd_sc_hd__a22o_1
X_14480_ _08348_ _08352_ _08353_ vssd1 vssd1 vccd1 vccd1 _08354_ sky130_fd_sc_hd__nand3_1
XFILLER_0_177_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11692_ game.CPU.applesa.ab.check_walls.above.walls\[62\] net256 _05580_ vssd1 vssd1
+ vccd1 vccd1 _05581_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_194_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ net681 _06965_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__or2_1
X_10643_ _04616_ _04689_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__or2_4
XANTENNA__17948__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12157__A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_341_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_354_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_311_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19345__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16150_ _02039_ _02044_ _02118_ _02161_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__o211a_1
X_13362_ _06677_ _06684_ net683 vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10574_ _03253_ net234 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__nor2_1
XANTENNA__10596__A1 game.CPU.applesa.ab.absxs.body_x\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_279_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15101_ net1203 net1229 game.CPU.applesa.ab.check_walls.above.walls\[129\] vssd1
+ vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__and3_1
XANTENNA__10596__B2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_341_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12313_ _06069_ _06070_ _06071_ _06163_ _06198_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__o311a_1
X_16081_ _03456_ net269 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13293_ net215 _07166_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__and2_1
XANTENNA__16720__A1 _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_267_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15032_ net1222 net1250 net817 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__and3_1
X_12244_ game.CPU.applesa.ab.check_walls.above.walls\[181\] net549 vssd1 vssd1 vccd1
+ vccd1 _06130_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_210_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19495__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19840_ clknet_leaf_36_clk game.writer.tracker.next_frame\[435\] net1351 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[435\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_310_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17276__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_283_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12175_ net806 net387 _06059_ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__a211o_1
XFILLER_0_294_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11126_ _03283_ net321 vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__xnor2_1
X_19771_ clknet_leaf_29_clk game.writer.tracker.next_frame\[366\] net1285 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[366\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15915__B net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16983_ _02461_ net90 _02666_ net1896 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[327\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16299__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17028__A2 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18722_ clknet_leaf_63_clk _01139_ _00459_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[96\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_147_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_322_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ _03252_ net406 net542 game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1
+ vccd1 vccd1 _04947_ sky130_fd_sc_hd__a22o_1
X_15934_ game.CPU.applesa.ab.check_walls.above.walls\[121\] net471 vssd1 vssd1 vccd1
+ vccd1 _01946_ sky130_fd_sc_hd__nor2_1
X_10008_ _04211_ _04214_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__and2_1
X_18653_ clknet_leaf_51_clk _01070_ _00390_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output49_A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16787__A1 _02465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15865_ _03323_ net337 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16787__B2 game.writer.tracker.frame\[200\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17604_ net2035 _03003_ _03018_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__o21ba_1
XANTENNA__15931__A game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14816_ game.CPU.randy.counter1.count\[14\] game.CPU.randy.counter1.count\[13\] _08621_
+ vssd1 vssd1 vccd1 vccd1 _08624_ sky130_fd_sc_hd__and3_1
X_18584_ clknet_leaf_12_clk _01004_ _00321_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[49\]
+ sky130_fd_sc_hd__dfrtp_4
X_15796_ game.CPU.applesa.ab.absxs.body_x\[50\] net467 net452 game.CPU.applesa.ab.absxs.body_y\[48\]
+ _01807_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14262__A2 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17535_ _02912_ _02915_ _02910_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_318_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_294_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11959_ net750 _05197_ _05846_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__a21oi_1
X_14747_ _08571_ _08572_ net55 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__and3b_1
XANTENNA__16539__B2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_236_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_317_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17200__A2 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17466_ _02887_ _02888_ _02890_ _02891_ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__o211a_1
X_14678_ game.CPU.randy.counter1.count1\[2\] _04352_ _08515_ _08516_ vssd1 vssd1 vccd1
+ vccd1 _08517_ sky130_fd_sc_hd__o211a_1
XFILLER_0_190_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19205_ clknet_leaf_70_clk _00018_ _00853_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.XMAX\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_333_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13629_ _07495_ _07502_ net278 vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__mux2_1
X_16417_ game.writer.tracker.frame\[44\] _02380_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_158_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19655__RESET_B net1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_317_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_251_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12067__A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17397_ game.CPU.kyle.L1.nextState\[3\] game.CPU.kyle.L1.nextState\[2\] vssd1 vssd1
+ vccd1 vccd1 _02827_ sky130_fd_sc_hd__nor2_2
XFILLER_0_305_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_305_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_307_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19136_ net1184 _00178_ _00807_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[181\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12576__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16348_ net195 _02334_ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__nand2_2
XANTENNA__14970__B1 net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18712__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19838__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16279_ net1008 _08400_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__nand2_1
X_19067_ net1185 _00102_ _00738_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[112\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13525__B2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18018_ net668 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
XANTENNA__09376__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_247_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout106 net110 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__buf_2
XANTENNA__16475__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout117 net118 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_4
XANTENNA__18862__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19988__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout128 net129 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_346_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19969_ clknet_leaf_42_clk game.writer.tracker.next_frame\[564\] net1326 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[564\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13289__B1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout139 _08601_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_169_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19581__Q game.writer.tracker.frame\[176\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14486__C1 _08184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13828__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ _03960_ _03961_ _03962_ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__a211o_1
XANTENNA__09823__B game.CPU.applesa.ab.absxs.body_x\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10969__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09901__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ net1082 game.CPU.applesa.ab.check_walls.above.walls\[171\] vssd1 vssd1 vccd1
+ vccd1 _03896_ sky130_fd_sc_hd__xor2_1
XANTENNA__16778__A1 _02450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19218__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09584_ net1150 game.CPU.applesa.ab.check_walls.above.walls\[21\] vssd1 vssd1 vccd1
+ vccd1 _03827_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_336_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13461__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14457__A game.CPU.applesa.ab.absxs.body_x\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout158_X net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_258_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1279_A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19368__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_271_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14005__A2 game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout704_A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19396__RESET_B net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10049__X _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1067_X net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13764__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12567__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16391__B _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12972__C1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18660__Q game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12264__X _06150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_347_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13516__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09018_ game.CPU.applesa.ab.absxs.body_x\[73\] vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__inv_2
X_10290_ net851 game.CPU.applesa.ab.x_final\[3\] game.CPU.applesa.ab.good_spot_next
+ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_269_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold160 game.writer.tracker.frame\[460\] vssd1 vssd1 vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17258__A2 _02300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold171 game.writer.tracker.frame\[324\] vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 game.writer.tracker.frame\[304\] vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16466__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 game.writer.tracker.frame\[215\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10750__A1 game.CPU.applesa.ab.absxs.body_y\[113\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_298_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout959_X net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 net651 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_4
Xfanout651 _08799_ vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13375__S0 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout662 net667 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_4
XANTENNA__09733__B game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13980_ net952 net828 vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__nand2_1
Xfanout673 net675 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_4
XFILLER_0_217_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout684 net685 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_2
XFILLER_0_260_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout695 net707 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_4
X_12931_ net511 _06804_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__or2_1
XANTENNA__16769__A1 _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10502__A1 game.CPU.applesa.ab.absxs.body_x\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_272_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16847__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10502__B2 game.CPU.applesa.ab.absxs.body_x\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_358_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13823__X _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15751__A game.CPU.applesa.ab.check_walls.above.walls\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_358_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ game.writer.tracker.frame\[258\] game.writer.tracker.frame\[259\] net997
+ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__mux2_1
X_15650_ _01655_ _01656_ _01660_ _01661_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__or4b_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16566__B _02415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_240_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14601_ _08458_ net741 _08457_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[4\]
+ sky130_fd_sc_hd__and3b_1
X_11813_ game.CPU.applesa.ab.check_walls.above.walls\[30\] net302 _05700_ vssd1 vssd1
+ vccd1 vccd1 _05701_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_205_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ game.CPU.applesa.ab.check_walls.above.walls\[89\] net474 vssd1 vssd1 vccd1
+ vccd1 _01593_ sky130_fd_sc_hd__xnor2_1
X_12793_ _06663_ _06664_ net687 vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__mux2_1
X_17320_ net2048 net732 _02762_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[568\]
+ sky130_fd_sc_hd__and3_1
X_14532_ _08401_ _08402_ _08405_ _08398_ _08397_ vssd1 vssd1 vccd1 vccd1 _08406_ sky130_fd_sc_hd__a32o_1
X_11744_ game.CPU.applesa.ab.check_walls.above.walls\[156\] net390 net299 game.CPU.applesa.ab.check_walls.above.walls\[158\]
+ _05629_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__a221o_1
XANTENNA__10805__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13204__A0 game.writer.tracker.frame\[432\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17251_ net70 _02368_ _02743_ net1924 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[518\]
+ sky130_fd_sc_hd__a2bb2o_1
X_14463_ game.CPU.applesa.ab.absxs.body_y\[61\] net965 vssd1 vssd1 vccd1 vccd1 _08337_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__18735__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11503__B net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11675_ game.CPU.applesa.ab.check_walls.above.walls\[124\] net249 _05561_ _05562_
+ _05563_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__o2111a_1
XANTENNA__16582__A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16941__A1 _02382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13414_ net287 _07278_ _07287_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__a21oi_1
X_16202_ game.CPU.applesa.ab.check_walls.above.walls\[11\] net463 net447 net830 _01686_
+ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__a221o_1
XANTENNA__12558__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12318__C _06201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17182_ _02485_ net74 _02726_ net1524 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[466\]
+ sky130_fd_sc_hd__a22o_1
X_10626_ _03240_ net327 vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__nor2_1
X_14394_ game.CPU.applesa.ab.absxs.body_x\[69\] net1067 vssd1 vssd1 vccd1 vccd1 _08268_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_180_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16133_ game.CPU.applesa.ab.absxs.body_x\[23\] net460 net440 game.CPU.applesa.ab.absxs.body_y\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__a2bb2o_1
X_13345_ net488 _06612_ _07218_ net686 vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10834__S _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10557_ net754 _04644_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__nor2_4
XFILLER_0_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13210__S net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18885__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16064_ game.CPU.applesa.ab.check_walls.above.walls\[194\] net466 vssd1 vssd1 vccd1
+ vccd1 _02076_ sky130_fd_sc_hd__nor2_1
X_13276_ _07148_ _07149_ net476 vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_310_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10488_ game.CPU.applesa.ab.absxs.body_x\[84\] _04610_ _04611_ game.CPU.applesa.ab.absxs.body_x\[80\]
+ vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_324_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15015_ net1221 net1249 game.CPU.applesa.ab.check_walls.above.walls\[43\] vssd1 vssd1
+ vccd1 vccd1 _00234_ sky130_fd_sc_hd__and3_1
XANTENNA__17249__A2 _02454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12227_ net809 net417 _06112_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_248_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16457__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19823_ clknet_leaf_39_clk game.writer.tracker.next_frame\[418\] net1350 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[418\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15645__B net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ _05254_ _05255_ _05257_ _05259_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__or4b_1
XANTENNA__10741__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ _03276_ net323 vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__xnor2_1
X_19754_ clknet_leaf_25_clk game.writer.tracker.next_frame\[349\] net1321 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[349\] sky130_fd_sc_hd__dfrtp_1
X_16966_ _02428_ net94 _02660_ net1746 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[316\]
+ sky130_fd_sc_hd__a22o_1
X_12089_ net828 net292 vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__xor2_1
XFILLER_0_251_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11549__A1_N game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18705_ clknet_leaf_31_clk _01122_ _00442_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[59\]
+ sky130_fd_sc_hd__dfrtp_2
X_15917_ _03449_ net449 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__nand2_1
X_19685_ clknet_leaf_34_clk game.writer.tracker.next_frame\[280\] net1322 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[280\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13691__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16897_ net145 _02291_ net86 net714 vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_242_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18636_ clknet_leaf_64_clk _01053_ _00373_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_204_Left_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15848_ game.CPU.applesa.ab.absxs.body_x\[79\] net460 net339 _03301_ vssd1 vssd1
+ vccd1 vccd1 _01860_ sky130_fd_sc_hd__o22a_1
XANTENNA__19510__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18745__Q game.CPU.applesa.ab.absxs.body_x\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_91_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18567_ clknet_leaf_9_clk _00987_ _00304_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_15779_ game.CPU.applesa.ab.absxs.body_x\[104\] net355 net344 _03252_ vssd1 vssd1
+ vccd1 vccd1 _01791_ sky130_fd_sc_hd__a22o_1
XFILLER_0_332_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17518_ net1259 game.CPU.speed1.Qa\[1\] net427 _02937_ net1243 vssd1 vssd1 vccd1
+ vccd1 _02946_ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17185__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_50_clk_X clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18498_ net584 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__inv_2
XANTENNA__12509__B net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11413__B net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17449_ _02872_ _02874_ _02877_ _08808_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__o31ai_4
XANTENNA__19660__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16932__A1 _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19119_ net1182 _00159_ _00790_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[164\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_213_Left_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_65_clk_X clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12525__A game.CPU.applesa.ab.absxs.body_x\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_298_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16160__A2 _02167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12244__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_246_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10045__A net1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09834__A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16999__A1 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_226_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19040__CLK net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10732__A1 game.CPU.applesa.ab.absxs.body_y\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_342_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18608__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14474__A2 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ net894 net817 _03416_ net1131 _03947_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_222_Left_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09886__C1 _03608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09636_ _03869_ _03870_ _03877_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__a22o_1
XANTENNA__19190__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18655__Q game.CPU.applesa.ab.absxs.body_y\[69\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_328_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18758__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ net1126 _03299_ game.CPU.applesa.ab.absxs.body_y\[76\] net891 _03807_ vssd1
+ vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_242_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19577__RESET_B net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1184_X net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout919_A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11604__A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_clk_X clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17176__A1 _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09498_ net1095 _03407_ _03409_ net1151 _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__a221o_1
XANTENNA__10799__A1 game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10799__B2 game.CPU.applesa.ab.absxs.body_y\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11996__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1351_X net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11460_ game.CPU.applesa.ab.check_walls.above.walls\[21\] net317 vssd1 vssd1 vccd1
+ vccd1 _05349_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_231_Left_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19486__Q game.writer.tracker.frame\[81\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_clk_X clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11748__B1 _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10411_ net1260 _04556_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__or2_1
XFILLER_0_351_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ net805 net257 vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_277_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13130_ game.writer.tracker.frame\[130\] game.writer.tracker.frame\[131\] net1005
+ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_289_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10342_ net1720 _04506_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13061_ game.writer.tracker.frame\[248\] game.writer.tracker.frame\[249\] net1031
+ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__mux2_1
XANTENNA__15746__A game.CPU.applesa.ab.check_walls.above.walls\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10273_ net1170 _04362_ _04367_ net1171 _04465_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout90_X net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_249_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12012_ _05895_ _05896_ _05897_ _05898_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_280_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11993__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17100__A1 _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16820_ net156 _02359_ net98 net715 vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__o31a_1
XANTENNA__17961__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_306_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09463__B net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout470 _08420_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19533__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout481 net483 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15662__B2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout492 net493 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_260_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16751_ net164 net67 net101 _02585_ net1511 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[175\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__11901__A2_N net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13963_ _07833_ _07834_ _07836_ _07832_ vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__a211o_1
XANTENNA__09877__C1 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09341__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15702_ game.CPU.applesa.ab.check_walls.above.walls\[156\] net342 vssd1 vssd1 vccd1
+ vccd1 _01714_ sky130_fd_sc_hd__nand2_1
XANTENNA__09341__B2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19470_ clknet_leaf_35_clk game.writer.tracker.next_frame\[65\] net1345 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[65\] sky130_fd_sc_hd__dfrtp_2
X_12914_ net211 _06785_ _06787_ net277 vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__a31o_1
X_16682_ net1992 _02554_ net62 _02452_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[131\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13894_ net873 game.CPU.applesa.ab.check_walls.above.walls\[59\] game.CPU.applesa.ab.check_walls.above.walls\[61\]
+ net864 _07767_ vssd1 vssd1 vccd1 vccd1 _07768_ sky130_fd_sc_hd__a221o_1
XFILLER_0_201_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_204_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18421_ net626 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__inv_2
X_12845_ game.writer.tracker.frame\[308\] game.writer.tracker.frame\[309\] net1028
+ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__mux2_1
X_15633_ _01640_ _01642_ _01643_ _01644_ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__or4_1
XANTENNA__19683__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14097__A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11514__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_291_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ net593 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__inv_2
XANTENNA__13976__A1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12776_ game.writer.tracker.frame\[124\] game.writer.tracker.frame\[125\] net1033
+ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__mux2_1
XANTENNA__17167__A1 _02461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15564_ _08937_ _01581_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13976__B2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17303_ net1943 net723 _02757_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[556\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_185_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11233__B net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14515_ _03206_ net1060 net958 _03205_ _08386_ vssd1 vssd1 vccd1 vccd1 _08389_ sky130_fd_sc_hd__a221o_1
X_11727_ game.CPU.applesa.ab.check_walls.above.walls\[76\] net395 net307 net813 vssd1
+ vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_138_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15495_ net676 _01506_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18283_ net622 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XANTENNA__16914__A1 _02491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09329__A1_N net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11801__X _05689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17234_ net154 _02422_ net79 _02739_ net2049 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[505\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_315_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_299_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14446_ _08314_ _08315_ _08316_ _08317_ vssd1 vssd1 vccd1 vccd1 _08320_ sky130_fd_sc_hd__a22o_1
X_11658_ game.CPU.applesa.ab.check_walls.above.walls\[14\] net256 net317 net830 vssd1
+ vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09197__Y _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10609_ game.CPU.applesa.ab.absxs.body_x\[82\] _04673_ _04674_ game.CPU.applesa.ab.absxs.body_x\[78\]
+ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17165_ _02458_ net78 _02722_ net1977 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[453\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14377_ game.CPU.applesa.ab.absxs.body_x\[83\] net1044 vssd1 vssd1 vccd1 vccd1 _08251_
+ sky130_fd_sc_hd__xnor2_1
X_11589_ game.CPU.applesa.ab.check_walls.above.walls\[106\] net767 vssd1 vssd1 vccd1
+ vccd1 _05478_ sky130_fd_sc_hd__xor2_2
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13328_ net200 _07201_ net276 vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__a21o_1
X_16116_ game.CPU.applesa.ab.absxs.body_x\[69\] net473 vssd1 vssd1 vccd1 vccd1 _02128_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17096_ _02491_ net60 _02700_ net1610 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[406\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16142__A2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19063__CLK net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_310_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15656__A game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13259_ game.writer.tracker.frame\[450\] game.writer.tracker.frame\[451\] net1014
+ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_268_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16047_ _02049_ _02056_ _02057_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__or3_1
XANTENNA__12703__A2 _06571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_244_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11911__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19806_ clknet_leaf_38_clk game.writer.tracker.next_frame\[401\] net1328 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[401\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_257_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17998_ net637 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__inv_2
XFILLER_0_223_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19737_ clknet_leaf_18_clk game.writer.tracker.next_frame\[332\] net1289 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[332\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_193_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16949_ net163 net67 net87 _02656_ net1555 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[303\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__11408__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16487__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18900__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09332__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13904__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09332__B2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19668_ clknet_leaf_29_clk game.writer.tracker.next_frame\[263\] net1285 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[263\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_343_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14208__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09883__A2 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09421_ net915 game.CPU.applesa.ab.absxs.body_x\[97\] game.CPU.applesa.ab.absxs.body_x\[96\]
+ net911 _03662_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__a221o_1
X_18619_ clknet_leaf_13_clk _01036_ _00356_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[113\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_189_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19599_ clknet_leaf_22_clk game.writer.tracker.next_frame\[194\] net1343 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[194\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19670__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ net917 game.CPU.applesa.ab.absxs.body_x\[9\] game.CPU.applesa.ab.absxs.body_y\[9\]
+ net899 _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_47_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13967__A1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_255_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13967__B2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12239__B net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11143__B net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09283_ game.CPU.applesa.ab.check_walls.above.walls\[192\] game.CPU.applesa.ab.check_walls.above.walls\[193\]
+ game.CPU.applesa.ab.check_walls.above.walls\[194\] game.CPU.applesa.ab.check_walls.above.walls\[195\]
+ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__nor4_1
XANTENNA__11442__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12954__S net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_30_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10982__B net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19406__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12255__A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14392__B2 game.CPU.applesa.ab.absxs.body_y\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout402_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17330__A1 _01454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_344_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_45_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1311_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_266_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19556__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09564__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10705__A1 game.CPU.applesa.ab.absxs.body_y\[69\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12702__B _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17094__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__A1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A _03374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16323__C_N _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08998_ game.CPU.applesa.ab.absxs.body_x\[31\] vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__inv_2
XANTENNA__14447__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_317_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11318__B _05206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18580__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12631__A2_N net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13750__S0 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ _03288_ net325 vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_253_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_355_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09619_ net1094 game.CPU.applesa.ab.check_walls.above.walls\[2\] vssd1 vssd1 vccd1
+ vccd1 _03862_ sky130_fd_sc_hd__xor2_1
X_10891_ _04448_ _04455_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__nand2_1
XANTENNA__10649__S _04690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13025__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_119_Left_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_329_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_277_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12630_ _06352_ _06468_ _06505_ _06506_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__or4_4
XANTENNA__10876__C game.CPU.applesa.ab.apple_possible\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11334__A game.CPU.applesa.ab.check_walls.above.walls\[83\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17149__A1 _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_356_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11053__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12561_ _06437_ _06429_ _06431_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__or3b_2
XANTENNA__12864__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14300_ game.CPU.applesa.ab.absxs.body_x\[30\] net1054 vssd1 vssd1 vccd1 vccd1 _08174_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11512_ net777 _05400_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_309_Left_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09739__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15280_ _01264_ _08830_ _08833_ vssd1 vssd1 vccd1 vccd1 _08834_ sky130_fd_sc_hd__a21oi_1
X_12492_ game.CPU.applesa.ab.absxs.body_x\[82\] net370 vssd1 vssd1 vccd1 vccd1 _06369_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10892__B net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12918__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14231_ _08094_ _08095_ _08096_ _08104_ vssd1 vssd1 vccd1 vccd1 _08105_ sky130_fd_sc_hd__or4_1
XFILLER_0_297_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11443_ game.CPU.applesa.ab.check_walls.above.walls\[74\] net768 vssd1 vssd1 vccd1
+ vccd1 _05332_ sky130_fd_sc_hd__xor2_2
XFILLER_0_123_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12165__A game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire178 net179 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_2
X_14162_ net1112 net1075 vssd1 vssd1 vccd1 vccd1 _08036_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11374_ net822 _05207_ _05262_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__o21ba_1
XANTENNA__16124__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17321__B2 _02275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_308_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13113_ net482 _06986_ net676 vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__a21o_1
XANTENNA__14135__A1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Left_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15588__A2_N net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13569__S0 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10325_ net740 _04493_ net1910 vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_265_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18970_ net1200 _00154_ _00641_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14093_ net885 game.CPU.applesa.ab.check_walls.above.walls\[9\] game.CPU.applesa.ab.check_walls.above.walls\[12\]
+ net870 _07966_ vssd1 vssd1 vccd1 vccd1 _07967_ sky130_fd_sc_hd__a221o_1
XANTENNA__14135__B2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12146__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13044_ _06916_ _06917_ net504 vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__mux2_1
X_17921_ net605 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__inv_2
X_10256_ net1173 _04446_ _04448_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13894__B1 game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1210 net1216 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__buf_2
XANTENNA__09562__A1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18923__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1221 game.CPU.walls.rand_wall.start_enable vssd1 vssd1 vccd1 vccd1 net1221
+ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_318_Left_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17852_ _03172_ _03176_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__nor2_1
XANTENNA__09562__B2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1232 net1257 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__clkbuf_2
X_10187_ _04372_ _04379_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1243 net1257 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__clkbuf_4
Xfanout1254 net1255 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__clkbuf_2
X_16803_ net150 _02327_ net104 _02601_ net1866 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[212\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_273_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1265 game.CPU.applesa.ab.absxs.body_x\[103\] vssd1 vssd1 vccd1 vccd1 net1265
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11228__B net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1276 net1277 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13646__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1287 net1288 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15923__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17783_ _03128_ _03129_ _03131_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__and3_1
X_14995_ net1228 net1252 game.CPU.applesa.ab.check_walls.above.walls\[23\] vssd1 vssd1
+ vccd1 vccd1 _00212_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_58_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_8
Xfanout1298 net1300 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__clkbuf_4
X_19522_ clknet_leaf_21_clk game.writer.tracker.next_frame\[117\] net1335 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[117\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13741__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16734_ net184 _02521_ net101 _02580_ net1552 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[164\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_31_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13946_ net993 _03418_ _03420_ net956 _07816_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_137_Left_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output31_A net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_319_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19453_ clknet_leaf_43_clk game.writer.tracker.next_frame\[48\] net1327 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[48\] sky130_fd_sc_hd__dfrtp_1
X_16665_ _02243_ net157 _02432_ net731 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__o31a_1
X_13877_ net1070 _03436_ game.CPU.applesa.ab.check_walls.above.walls\[110\] net852
+ vssd1 vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__o22a_1
XFILLER_0_186_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18404_ net602 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__inv_2
X_15616_ game.CPU.applesa.ab.check_walls.above.walls\[86\] net333 vssd1 vssd1 vccd1
+ vccd1 _01628_ sky130_fd_sc_hd__nand2_1
X_12828_ _06634_ _06636_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__xnor2_2
X_19384_ clknet_leaf_3_clk _01390_ _00964_ vssd1 vssd1 vccd1 vccd1 game.CPU.bodymain1.main.score\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_335_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16596_ net129 net56 _02439_ _02510_ net2045 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[96\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_201_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12059__B net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_347_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19429__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18335_ net592 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_327_Left_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15547_ _06551_ _06556_ _01473_ _01533_ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_328_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12759_ _06551_ _06555_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__and2_2
XFILLER_0_173_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14555__A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18266_ net622 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
X_15478_ _01456_ _01463_ _01499_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12909__C1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17217_ net53 net142 net119 _02735_ net1497 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[492\]
+ sky130_fd_sc_hd__a32o_1
X_14429_ game.CPU.applesa.ab.absxs.body_y\[26\] net949 vssd1 vssd1 vccd1 vccd1 _08303_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09368__B game.CPU.applesa.ab.check_walls.above.walls\[32\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16770__A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_287_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18197_ net581 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__inv_2
XANTENNA__15089__C net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_250_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19579__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17148_ _02423_ net58 _02716_ net1484 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[442\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17312__A1 _02276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19854__Q game.writer.tracker.frame\[449\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14126__A1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_272_Right_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14126__B2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09970_ _04196_ _04197_ net1136 vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__o21a_1
X_17079_ _02466_ net57 _02696_ game.writer.tracker.frame\[393\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[393\] sky130_fd_sc_hd__a22o_1
XANTENNA__12137__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13334__C1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_336_Left_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12522__B net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_354_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13637__A0 game.writer.tracker.frame\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15833__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11138__B net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12949__S net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout185_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_211_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17379__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10977__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout352_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__A3 _04594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1094_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ _03641_ _03642_ _03644_ _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__or4b_1
X_20037__1385 vssd1 vssd1 vccd1 vccd1 net1385 _20037__1385/LO sky130_fd_sc_hd__conb_1
XANTENNA__10871__B1 game.CPU.randy.counter1.count\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_326_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09335_ net1128 game.CPU.applesa.ab.absxs.body_y\[91\] vssd1 vssd1 vccd1 vccd1 _03578_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12612__A1 game.CPU.applesa.ab.absxs.body_y\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_319_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10993__A game.CPU.applesa.ab.absxs.body_x\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_353_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout617_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17536__D1 _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17000__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_X net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1359_A net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_350_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09559__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ game.CPU.randy.counter1.count\[2\] vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__inv_2
XANTENNA__14184__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_279_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11601__B net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09197_ net794 vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__inv_2
XANTENNA__16680__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1147_X net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_214_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09993__S _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout986_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16657__A3 _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1314_X net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13325__C1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout98_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ net1629 _04312_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__or2_1
XFILLER_0_286_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11090_ game.CPU.applesa.ab.absxs.body_x\[60\] net324 vssd1 vssd1 vccd1 vccd1 _04980_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09544__A1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_186_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ net1171 _04218_ _04237_ net1170 _04248_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__a221o_1
XANTENNA__12774__S1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_328_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold20 game.CPU.walls.abc.number\[0\] vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 game.CPU.walls.abc.number\[5\] vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_303_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold42 game.CPU.applesa.normal1.number\[5\] vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15743__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11048__B net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold53 game.CPU.applesa.ab.absxs.body_x\[0\] vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 game.CPU.applesa.ab.absxs.body_x\[3\] vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout941_X net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold75 game.CPU.applesa.twoapples.count\[3\] vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ net514 _07669_ _07670_ _07673_ net230 vssd1 vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__a311o_1
Xhold86 game.writer.tracker.frame\[171\] vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09741__B game.CPU.applesa.ab.check_walls.above.walls\[66\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold97 game.CPU.clock1.counter\[10\] vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15462__C _01454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14780_ game.CPU.randy.counter1.count\[18\] _04486_ _08600_ vssd1 vssd1 vccd1 vccd1
+ _08601_ sky130_fd_sc_hd__nor3_1
X_11992_ net826 net553 vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout53_X net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14359__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13731_ game.writer.tracker.frame\[222\] net845 net837 game.writer.tracker.frame\[221\]
+ vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__o22a_1
X_10943_ _03315_ net543 vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__nand2_1
XANTENNA__19004__Q game.CPU.applesa.ab.check_walls.above.walls\[49\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_280_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_201_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16450_ net1820 _02406_ _02409_ net137 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[51\]
+ sky130_fd_sc_hd__a22o_1
X_13662_ game.writer.tracker.frame\[9\] game.writer.tracker.frame\[11\] game.writer.tracker.frame\[12\]
+ game.writer.tracker.frame\[10\] net970 net1002 vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__mux4_1
X_10874_ game.CPU.applesa.ab.apple_possible\[4\] net759 vssd1 vssd1 vccd1 vccd1 _04776_
+ sky130_fd_sc_hd__nand2_1
Xclkbuf_3_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_356_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15401_ game.writer.updater.commands.count\[13\] _01427_ _01428_ game.writer.updater.commands.count\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__a31o_1
XANTENNA__17022__Y _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12613_ _06425_ _06426_ _06427_ _06458_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__and4_1
X_13593_ game.writer.tracker.frame\[377\] game.writer.tracker.frame\[379\] game.writer.tracker.frame\[380\]
+ game.writer.tracker.frame\[378\] net979 net1032 vssd1 vssd1 vccd1 vccd1 _07467_
+ sky130_fd_sc_hd__mux4_1
X_16381_ _02314_ _02356_ _02358_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__o21ba_4
XTAP_TAPCELL_ROW_197_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_356_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18120_ net582 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_139_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_344_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_325_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15332_ game.CPU.applesa.twomode.number\[3\] _08871_ vssd1 vssd1 vccd1 vccd1 _08875_
+ sky130_fd_sc_hd__or2_1
X_12544_ game.CPU.applesa.ab.absxs.body_y\[43\] net367 vssd1 vssd1 vccd1 vccd1 _06421_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_314_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19721__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14094__B game.CPU.applesa.ab.check_walls.above.walls\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18051_ net659 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__inv_2
XANTENNA__11511__B net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12475_ game.CPU.applesa.ab.absxs.body_x\[57\] net379 vssd1 vssd1 vccd1 vccd1 _06352_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15263_ _08817_ _01262_ vssd1 vssd1 vccd1 vccd1 _08819_ sky130_fd_sc_hd__nor2_1
XFILLER_0_289_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17002_ _02327_ net83 _02672_ net2001 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[340\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13564__C1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14214_ _03229_ net1054 net949 _03296_ _08082_ vssd1 vssd1 vccd1 vccd1 _08088_ sky130_fd_sc_hd__a221o_1
X_11426_ net826 net252 vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15194_ game.CPU.applesa.normal1.counter_normal game.CPU.applesa.normal1.number\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08764_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _02179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_300_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15918__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_340_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09783__A1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14145_ _07847_ _07853_ _08018_ vssd1 vssd1 vccd1 vccd1 _08019_ sky130_fd_sc_hd__o21bai_2
XANTENNA__16648__A3 _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19871__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09783__B2 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ net791 net254 vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_78_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11590__B2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10308_ game.CPU.randy.f1.a1.count\[8\] game.CPU.randy.f1.a1.count\[7\] _04490_ vssd1
+ vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__and3_1
XFILLER_0_265_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18953_ clknet_leaf_67_clk net1416 _00624_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14076_ game.CPU.applesa.ab.YMAX\[1\] net862 game.CPU.applesa.ab.YMAX\[0\] net867
+ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__o211a_1
X_11288_ _04981_ _04985_ _05176_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__or4_4
XANTENNA__13867__B1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12342__B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17058__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _06863_ _06882_ net698 vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__mux2_1
X_17904_ net669 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__inv_2
XANTENNA__09535__A1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_265_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10239_ _04376_ _04378_ _04393_ _04430_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__o22a_1
XANTENNA__15934__A game.CPU.applesa.ab.check_walls.above.walls\[121\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09535__B2 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18884_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[14\] _00579_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_238_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11342__A1 _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1040 net1041 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11342__B2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1051 game.CPU.applesa.x\[3\] vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_8
X_17835_ game.writer.updater.commands.count\[6\] _03161_ vssd1 vssd1 vccd1 vccd1 _03164_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1062 game.CPU.applesa.x\[1\] vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_163_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15653__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1073 net1077 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__buf_2
Xfanout1084 net1088 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_145_Left_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13454__A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1095 game.CPU.applesa.ab.snake_head_x\[2\] vssd1 vssd1 vccd1 vccd1 net1095
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__16281__B2 _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09651__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16820__A3 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13095__A1 _06967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17766_ game.CPU.applesa.twoapples.count_luck\[4\] _03116_ game.CPU.applesa.twoapples.count_luck\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__a21o_1
X_14978_ net1225 net1252 game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1
+ vccd1 vccd1 _00143_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19505_ clknet_leaf_14_clk game.writer.tracker.next_frame\[100\] net1282 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[100\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_221_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16717_ net160 _02341_ net109 _02572_ net1638 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[154\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__13190__S1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19251__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13929_ net1063 game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1 vssd1 vccd1
+ vccd1 _07803_ sky130_fd_sc_hd__or2_1
X_17697_ game.CPU.walls.rand_wall.count\[0\] net1175 vssd1 vssd1 vccd1 vccd1 _03076_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_297_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19436_ clknet_leaf_41_clk game.writer.tracker.next_frame\[31\] net1332 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[31\] sky130_fd_sc_hd__dfrtp_1
X_16648_ net190 net125 _02410_ _02540_ net1622 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[116\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_239_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_347_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16484__B _02351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_252_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19367_ clknet_leaf_71_clk _01373_ _00948_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location2\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_335_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16579_ net118 _02499_ net558 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_341_Right_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_340_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09120_ net1065 vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__inv_2
XANTENNA__09379__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10605__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18318_ net615 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19298_ clknet_leaf_69_clk net319 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.x_final\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17533__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_154_Left_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12517__B net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09051_ game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__inv_2
XANTENNA__11421__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18249_ net644 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
XFILLER_0_199_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_331_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold501 game.writer.tracker.frame\[418\] vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15828__B net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10908__A1 game.CPU.applesa.enable_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold512 game.writer.tracker.frame\[221\] vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 game.writer.tracker.frame\[398\] vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09774__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_344_Left_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold534 game.writer.tracker.frame\[550\] vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09774__B2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold545 game.writer.tracker.frame\[192\] vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09826__B game.CPU.applesa.ab.absxs.body_y\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold556 game.writer.tracker.frame\[36\] vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold567 game.writer.tracker.frame\[119\] vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_268_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13307__C1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold578 game.writer.tracker.frame\[30\] vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 game.writer.tracker.frame\[185\] vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _04175_ _04184_ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__and2_1
XANTENNA__16499__X _02444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_263_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12252__B net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ _03876_ _03880_ _03941_ _04124_ _04126_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_209_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1107_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_163_Left_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12530__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout188_X net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout567_A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09829__A2 game.CPU.applesa.ab.absxs.body_y\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14283__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_353_Left_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_352_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout734_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_X net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19744__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16575__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_274_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_314_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_216_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13303__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_172_Left_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09318_ net1131 game.CPU.applesa.ab.absxs.body_y\[67\] vssd1 vssd1 vccd1 vccd1 _03561_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13794__C1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09289__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ game.CPU.applesa.ab.absxs.body_x\[109\] _04665_ _04666_ game.CPU.applesa.ab.absxs.body_x\[105\]
+ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_353_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16681__Y _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12427__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11331__B net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09249_ game.CPU.randy.counter1.count1\[16\] vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__inv_2
XANTENNA__19894__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12349__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13546__C1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09576__X _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_279_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ _05890_ _06145_ _05888_ _05889_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__or4bb_1
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15738__B net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout989_X net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ _03228_ net546 vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__nand2_1
X_12191_ game.CPU.applesa.ab.check_walls.above.walls\[127\] net422 vssd1 vssd1 vccd1
+ vccd1 _06077_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10515__X _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput10 net10 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XANTENNA__19124__CLK net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
X_11142_ _03262_ net326 vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__xnor2_1
Xoutput43 net43 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XANTENNA__13849__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_290_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_227_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_181_Left_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15950_ _01958_ _01959_ _01960_ _01961_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__or4_1
X_11073_ game.CPU.applesa.ab.absxs.body_x\[41\] net413 vssd1 vssd1 vccd1 vccd1 _04963_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_247_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19702__RESET_B net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ net1164 game.CPU.applesa.out_random_2\[2\] vssd1 vssd1 vccd1 vccd1 _04232_
+ sky130_fd_sc_hd__nand2_1
X_14901_ net1144 _08426_ vssd1 vssd1 vccd1 vccd1 _08678_ sky130_fd_sc_hd__nor2_1
X_15881_ _03452_ net346 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__nor2_1
XANTENNA__19274__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17620_ net2037 _03027_ net429 vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_355_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14832_ game.CPU.randy.f1.c1.count\[0\] game.CPU.randy.f1.c1.count\[1\] game.CPU.randy.f1.c1.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _08634_ sky130_fd_sc_hd__a21o_1
XFILLER_0_208_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14274__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14089__B game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _02783_ _02873_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__nor2_1
XANTENNA__11506__B net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14763_ game.CPU.randy.counter1.count\[12\] game.CPU.randy.counter1.count\[8\] net265
+ vssd1 vssd1 vccd1 vccd1 _08584_ sky130_fd_sc_hd__o21a_1
XANTENNA__11627__A2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11975_ game.CPU.applesa.ab.check_walls.above.walls\[150\] net288 vssd1 vssd1 vccd1
+ vccd1 _05862_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_291_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_316_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _02283_ net196 _02399_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__or3_1
XANTENNA__17212__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13714_ _07586_ _07587_ net477 vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10926_ net396 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.next_head\[7\] sky130_fd_sc_hd__inv_2
X_17482_ _02902_ _02904_ _02907_ _02909_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__o31ai_1
X_14694_ _08531_ _08532_ vssd1 vssd1 vccd1 vccd1 _08533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_357_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_224_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19221_ clknet_leaf_69_clk _01315_ _00860_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_location\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_16433_ net195 _02353_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__nor2_8
XANTENNA__18573__Q game.CPU.applesa.ab.absxs.body_y\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_345_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13645_ game.writer.tracker.frame\[25\] net838 net674 game.writer.tracker.frame\[28\]
+ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__o22a_1
X_10857_ game.CPU.randy.counter1.count\[16\] _03497_ _04740_ vssd1 vssd1 vccd1 vccd1
+ _04760_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12588__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13785__C1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19152_ net1187 _00195_ _00823_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[197\]
+ sky130_fd_sc_hd__dfrtp_4
X_16364_ net2054 net737 _02346_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[28\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_344_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13576_ game.writer.tracker.frame\[325\] game.writer.tracker.frame\[327\] game.writer.tracker.frame\[328\]
+ game.writer.tracker.frame\[326\] net978 net1027 vssd1 vssd1 vccd1 vccd1 _07450_
+ sky130_fd_sc_hd__mux4_1
X_10788_ net932 game.CPU.applesa.ab.absxs.body_y\[46\] net561 _04725_ vssd1 vssd1
+ vccd1 vccd1 _01005_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_344_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ net632 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__inv_2
XANTENNA__11241__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15315_ game.CPU.applesa.twomode.number\[0\] _08856_ vssd1 vssd1 vccd1 vccd1 _08861_
+ sky130_fd_sc_hd__or2_1
XANTENNA__15526__B1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15929__A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19083_ net1177 _00119_ _00754_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[128\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12527_ game.CPU.applesa.ab.absxs.body_y\[96\] net359 vssd1 vssd1 vccd1 vccd1 _06404_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16869__A3 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16295_ net1008 net866 _01516_ _02294_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a31o_1
XANTENNA__16133__A2_N net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18034_ net590 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__inv_2
X_15246_ game.CPU.kyle.L1.cnt_500hz\[7\] game.CPU.kyle.L1.cnt_500hz\[8\] game.CPU.kyle.L1.cnt_500hz\[10\]
+ game.CPU.kyle.L1.cnt_500hz\[11\] vssd1 vssd1 vccd1 vccd1 _08807_ sky130_fd_sc_hd__and4_1
X_12458_ _06328_ _06330_ _06332_ _06334_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__or4b_1
XFILLER_0_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15541__A3 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_313_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11012__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_327_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11409_ net799 net251 vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15177_ _04577_ _08752_ vssd1 vssd1 vccd1 vccd1 _08753_ sky130_fd_sc_hd__and2_1
X_12389_ game.CPU.applesa.ab.absxs.body_y\[27\] net364 vssd1 vssd1 vccd1 vccd1 _06266_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__12353__A game.CPU.applesa.ab.absxs.body_y\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10366__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14128_ net1049 _03393_ game.CPU.applesa.ab.check_walls.above.walls\[31\] net859
+ _07999_ vssd1 vssd1 vccd1 vccd1 _08002_ sky130_fd_sc_hd__o221a_1
X_19985_ clknet_leaf_45_clk _01409_ net1304 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_20036__1384 vssd1 vssd1 vccd1 vccd1 net1384 _20036__1384/LO sky130_fd_sc_hd__conb_1
XANTENNA__12072__B net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_249_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19617__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_287_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18936_ clknet_leaf_15_clk net557 net1282 vssd1 vssd1 vccd1 vccd1 game.CPU.reset_button1.sync1.Q
+ sky130_fd_sc_hd__dfrtp_1
X_14059_ net886 game.CPU.applesa.ab.check_walls.above.walls\[144\] game.CPU.applesa.ab.check_walls.above.walls\[146\]
+ net877 _07932_ vssd1 vssd1 vccd1 vccd1 _07933_ sky130_fd_sc_hd__a221o_1
XFILLER_0_253_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19443__RESET_B net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11315__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12512__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16479__B _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18867_ clknet_leaf_0_clk _01258_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11866__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13184__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11256__X _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_265_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17818_ _08886_ _03150_ _03151_ net182 net1899 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__a32o_1
X_18798_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[1\] _00535_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10601__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18641__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14265__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19767__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11079__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17749_ net1271 _04308_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_221_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_351_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16557__A2 _02481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_336_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19419_ clknet_leaf_48_clk game.writer.tracker.next_frame\[14\] net1301 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[14\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18791__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout148_A _02270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13123__S net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13961__A1_N net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11432__A game.CPU.applesa.ab.check_walls.above.walls\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_335_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12247__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09103_ game.CPU.applesa.ab.absxs.body_y\[19\] vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__inv_2
XFILLER_0_323_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11251__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12962__S net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10048__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout315_A _05213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19147__CLK net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1057_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ game.CPU.applesa.ab.absxs.body_x\[17\] vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__inv_2
XANTENNA__10990__B net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14462__B net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11056__A2_N net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_300_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold320 game.writer.tracker.frame\[169\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 game.writer.tracker.frame\[441\] vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold342 game.writer.tracker.frame\[148\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1224_A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 game.writer.tracker.frame\[71\] vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 game.CPU.walls.rand_wall.count_luck\[2\] vssd1 vssd1 vccd1 vccd1 net1749
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 game.writer.tracker.frame\[117\] vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17285__A3 _02434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19297__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout684_A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold386 game.writer.tracker.frame\[544\] vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout800 game.CPU.applesa.ab.check_walls.above.walls\[111\] vssd1 vssd1 vccd1 vccd1
+ net800 sky130_fd_sc_hd__clkbuf_4
Xhold397 game.writer.tracker.frame\[121\] vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout811 game.CPU.applesa.ab.check_walls.above.walls\[79\] vssd1 vssd1 vccd1 vccd1
+ net811 sky130_fd_sc_hd__clkbuf_4
X_09936_ net1123 net1124 vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__nand2_4
Xfanout822 game.CPU.applesa.ab.check_walls.above.walls\[38\] vssd1 vssd1 vccd1 vccd1
+ net822 sky130_fd_sc_hd__buf_4
Xfanout844 net845 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__buf_2
XFILLER_0_271_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout855 _03377_ vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_183_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout866 _03375_ vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_4
XANTENNA__17037__A3 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18658__Q game.CPU.applesa.ab.absxs.body_y\[76\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09867_ net1111 game.CPU.applesa.ab.absxs.body_x\[108\] vssd1 vssd1 vccd1 vccd1 _04110_
+ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout877 net880 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__buf_4
Xfanout888 net889 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16245__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout949_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout899 net900 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_300_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16796__A2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14256__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09798_ _04033_ _04034_ _04035_ _04036_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__and4_1
XFILLER_0_325_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_222_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11326__B net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11760_ game.CPU.applesa.ab.check_walls.above.walls\[181\] net307 vssd1 vssd1 vccd1
+ vccd1 _05648_ sky130_fd_sc_hd__or2_1
XFILLER_0_339_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10711_ _03339_ net425 vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_327_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ _03415_ _05194_ _05206_ _05578_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__o311a_1
XFILLER_0_138_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13430_ _06948_ _06964_ net693 vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_194_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10642_ _04606_ _04615_ net848 vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__a21o_2
XFILLER_0_326_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12157__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13361_ _06670_ _06672_ _06678_ _06671_ net702 net493 vssd1 vssd1 vccd1 vccd1 _07235_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_311_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11061__B net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ net936 net1265 net234 _04659_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__a31o_1
XANTENNA__15749__A game.CPU.applesa.ab.check_walls.above.walls\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15100_ net1203 net1231 game.CPU.applesa.ab.check_walls.above.walls\[128\] vssd1
+ vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09747__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ _06196_ _06197_ _06194_ _06195_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__a211o_1
X_13292_ _06767_ _06770_ _06774_ _06769_ net706 net495 vssd1 vssd1 vccd1 vccd1 _07166_
+ sky130_fd_sc_hd__mux4_1
X_16080_ game.CPU.applesa.ab.check_walls.above.walls\[149\] net444 vssd1 vssd1 vccd1
+ vccd1 _02092_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_310_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16720__A2 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15031_ net1228 net1256 game.CPU.applesa.ab.check_walls.above.walls\[59\] vssd1 vssd1
+ vccd1 vccd1 _00251_ sky130_fd_sc_hd__and3_1
X_12243_ game.CPU.applesa.ab.check_walls.above.walls\[183\] net423 vssd1 vssd1 vccd1
+ vccd1 _06129_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13534__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_322_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17964__A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12173__A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12174_ net806 net387 _06060_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__o21ai_1
XANTENNA__17276__A3 _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_259_Left_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11125_ game.CPU.applesa.ab.absxs.body_y\[16\] net534 vssd1 vssd1 vccd1 vccd1 _05015_
+ sky130_fd_sc_hd__nand2_1
X_19770_ clknet_leaf_28_clk game.writer.tracker.next_frame\[365\] net1287 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[365\] sky130_fd_sc_hd__dfrtp_1
X_16982_ _02462_ net89 net558 vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__a21oi_2
XANTENNA__18664__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16299__B _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18721_ clknet_leaf_69_clk _01138_ _00458_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_147_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11056_ game.CPU.applesa.ab.absxs.body_y\[106\] net539 net545 game.CPU.applesa.ab.absxs.body_x\[107\]
+ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__a2bb2o_1
X_15933_ _03444_ net350 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__nor2_1
XANTENNA__18568__Q game.CPU.applesa.ab.absxs.body_y\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_322_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_290_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_290_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_290_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_250_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10007_ _04214_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18652_ clknet_leaf_51_clk _01069_ _00389_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[62\]
+ sky130_fd_sc_hd__dfrtp_4
X_15864_ game.CPU.applesa.ab.absxs.body_y\[112\] net452 vssd1 vssd1 vccd1 vccd1 _01876_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_216_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16787__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17603_ game.CPU.kyle.L1.cnt_20ms\[6\] _03003_ _03008_ net577 vssd1 vssd1 vccd1 vccd1
+ _03018_ sky130_fd_sc_hd__a31o_1
XFILLER_0_235_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14815_ net1687 _08621_ _08623_ vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_231_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18583_ clknet_leaf_12_clk _01003_ _00320_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[48\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15931__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15995__B1 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15795_ game.CPU.applesa.ab.absxs.body_y\[49\] net446 net355 game.CPU.applesa.ab.absxs.body_x\[48\]
+ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_98_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17534_ net1476 net264 _02880_ _02961_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__a22o_1
X_14746_ game.CPU.randy.counter1.count1\[13\] game.CPU.randy.counter1.count1\[12\]
+ _08565_ game.CPU.randy.counter1.count1\[14\] vssd1 vssd1 vccd1 vccd1 _08572_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_294_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_268_Left_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11958_ net750 _05197_ _05202_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_318_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14547__B _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_345_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_357_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_236_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10909_ _03213_ _04381_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17465_ _02890_ _02891_ _02887_ _02888_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__a211oi_1
X_14677_ game.CPU.randy.counter1.count1\[2\] _04352_ game.CPU.randy.counter1.count1\[1\]
+ vssd1 vssd1 vccd1 vccd1 _08516_ sky130_fd_sc_hd__a21o_1
XFILLER_0_357_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11889_ _05771_ _05772_ _05773_ _05776_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__and4_1
XANTENNA__10390__A1_N net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19204_ clknet_leaf_71_clk _00017_ _00852_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.XMAX\[1\]
+ sky130_fd_sc_hd__dfstp_4
X_16416_ net115 _02299_ net164 _02380_ net1572 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[43\]
+ sky130_fd_sc_hd__a32o_1
X_13628_ _07498_ _07501_ net228 vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__mux2_1
XANTENNA__13222__A1 game.writer.tracker.frame\[393\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_317_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17396_ net1258 _03219_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12067__B net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10036__A1 game.CPU.applesa.ab.XMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_317_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19135_ net1183 _00177_ _00806_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[180\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10036__B2 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13773__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12782__S net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16347_ net866 _02246_ net235 _02333_ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__a31o_1
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15659__A game.CPU.applesa.ab.check_walls.above.walls\[48\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13559_ game.writer.tracker.frame\[98\] net841 net672 game.writer.tracker.frame\[100\]
+ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_171_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18035__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_298_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12981__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09657__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19066_ net1186 _00101_ _00737_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_16278_ net2039 net718 _02281_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[7\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__16172__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14282__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18017_ net660 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__inv_2
XFILLER_0_313_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15229_ game.CPU.applesa.normal1.number\[6\] _08788_ vssd1 vssd1 vccd1 vccd1 _08793_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09376__B game.CPU.applesa.ab.check_walls.above.walls\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12083__A game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_277_Left_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15097__C net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16087__A2_N net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_247_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout107 net108 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13466__X _07340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16475__A1 _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout118 _02242_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__buf_4
XANTENNA__13907__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout129 _02344_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_4
X_19968_ clknet_leaf_42_clk game.writer.tracker.next_frame\[563\] net1330 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[563\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_253_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14486__B1 _08345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_253_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09721_ net1090 _03232_ _03298_ net1154 _03963_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__a221o_1
X_18919_ clknet_leaf_4_clk net1402 _00603_ vssd1 vssd1 vccd1 vccd1 game.CPU.down_button.eD1.Q2
+ sky130_fd_sc_hd__dfrtp_1
X_19899_ clknet_leaf_15_clk game.writer.tracker.next_frame\[494\] net1288 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[494\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11427__A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ net1154 net785 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__nand2_1
XANTENNA__16778__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10511__A2 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16496__Y _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11146__B net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15841__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09583_ net1140 net828 vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__xor2_1
XANTENNA__10050__B _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_286_Left_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09466__A2_N net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17114__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14457__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_258_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_309_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_271_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout432_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__A game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_336_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16950__A2 _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout220_X net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1341_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11775__A1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16163__B1 _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_295_Left_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_347_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09017_ game.CPU.applesa.ab.absxs.body_x\[80\] vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout899_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10506__A _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1227_X net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_269_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold150 game.CPU.applesa.ab.count_luck\[2\] vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09854__X _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19932__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 game.writer.tracker.frame\[476\] vssd1 vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 game.writer.tracker.frame\[380\] vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16466__A1 _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold183 game.writer.tracker.frame\[290\] vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13376__X _07250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 game.writer.tracker.frame\[139\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_245_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12721__A _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout80_A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_224_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14477__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 net632 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__buf_4
XANTENNA__10750__A2 _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_298_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout641 net642 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_4
Xfanout652 net655 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_4
X_09919_ net1084 _04155_ _04160_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__o21a_1
XANTENNA__13375__S1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout663 net667 vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__buf_4
Xfanout674 net675 vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12440__B net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout685 net692 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13028__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11337__A game.CPU.applesa.ab.check_walls.above.walls\[82\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12930_ _06709_ _06711_ net688 vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_272_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20039_ net1363 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
Xfanout696 net699 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_3_1_0_clk_X clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16769__A2 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11563__A2_N net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10502__A2 _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16847__B _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_272_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_358_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ game.writer.tracker.frame\[260\] game.writer.tracker.frame\[261\] net997
+ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15751__B net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_358_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14600_ game.CPU.clock1.counter\[3\] game.CPU.clock1.counter\[4\] _08455_ vssd1 vssd1
+ vccd1 vccd1 _08458_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_17_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ net826 net393 net302 game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1
+ vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__o22a_1
XFILLER_0_197_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15580_ game.CPU.applesa.ab.check_walls.above.walls\[95\] net433 vssd1 vssd1 vccd1
+ vccd1 _01592_ sky130_fd_sc_hd__xnor2_1
X_12792_ _06662_ _06665_ net688 vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__mux2_1
XANTENNA__13452__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14367__B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10895__B _04796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14531_ _07400_ _08403_ _07742_ vssd1 vssd1 vccd1 vccd1 _08405_ sky130_fd_sc_hd__a21o_1
XFILLER_0_185_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11743_ game.CPU.applesa.ab.check_walls.above.walls\[157\] net305 vssd1 vssd1 vccd1
+ vccd1 _05631_ sky130_fd_sc_hd__nand2_1
XANTENNA__17959__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17194__A2 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20035__1383 vssd1 vssd1 vccd1 vccd1 net1383 _20035__1383/LO sky130_fd_sc_hd__conb_1
XFILLER_0_83_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17250_ _02267_ _02275_ _02743_ net1824 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[517\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14462_ game.CPU.applesa.ab.absxs.body_x\[63\] net1048 vssd1 vssd1 vccd1 vccd1 _08336_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__14401__B1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11674_ net795 net314 vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16941__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16582__B _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13698__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16201_ _01921_ _02212_ _01922_ _02123_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__or4b_2
XFILLER_0_193_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13413_ net275 _07282_ _07286_ net243 vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__a31o_1
X_17181_ _02483_ net73 _02726_ net1650 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[465\]
+ sky130_fd_sc_hd__a22o_1
X_10625_ game.CPU.applesa.ab.absxs.body_x\[64\] _04679_ _04680_ game.CPU.applesa.ab.absxs.body_x\[60\]
+ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__a22o_1
XANTENNA__12318__D _06203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14393_ _08263_ _08265_ _08266_ vssd1 vssd1 vccd1 vccd1 _08267_ sky130_fd_sc_hd__or3_1
XANTENNA__11766__A1 game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09477__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16132_ game.CPU.applesa.ab.absxs.body_x\[23\] net460 net454 game.CPU.applesa.ab.absxs.body_y\[20\]
+ _02139_ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13344_ net511 _06762_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__or2_1
X_10556_ game.CPU.applesa.ab.absxs.body_x\[28\] net330 _04651_ net930 vssd1 vssd1
+ vccd1 vccd1 _01163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16063_ _03485_ net347 vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_297_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13275_ game.writer.tracker.frame\[490\] game.writer.tracker.frame\[491\] net995
+ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ game.CPU.applesa.ab.absxs.body_x\[85\] _04610_ _04611_ game.CPU.applesa.ab.absxs.body_x\[81\]
+ vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__a22o_1
X_15014_ net1220 net1248 game.CPU.applesa.ab.check_walls.above.walls\[42\] vssd1 vssd1
+ vccd1 vccd1 _00233_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_324_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12226_ _03425_ net547 vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16457__A1 _02234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_184_Right_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19822_ clknet_leaf_39_clk game.writer.tracker.next_frame\[417\] net1350 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[417\] sky130_fd_sc_hd__dfrtp_1
X_12157_ net824 net553 vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__or2_1
XFILLER_0_236_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_235_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14468__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10741__A2 game.CPU.applesa.ab.absxs.body_y\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_275_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11108_ _03277_ net416 vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__nand2_1
X_16965_ _02424_ net94 _02660_ net1783 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[315\]
+ sky130_fd_sc_hd__a22o_1
X_19753_ clknet_leaf_25_clk game.writer.tracker.next_frame\[348\] net1321 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[348\] sky130_fd_sc_hd__dfrtp_1
X_12088_ net827 net297 vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_263_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13140__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18704_ clknet_leaf_31_clk _01121_ _00441_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[58\]
+ sky130_fd_sc_hd__dfrtp_4
X_11039_ _04918_ _04919_ _04920_ _04921_ _04924_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a221o_1
X_15916_ net792 net336 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__or2_1
X_19684_ clknet_leaf_34_clk game.writer.tracker.next_frame\[279\] net1322 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[279\] sky130_fd_sc_hd__dfrtp_1
X_16896_ _02467_ net93 _02640_ net1717 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[266\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_246_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09895__B1 _03903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_242_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18635_ clknet_leaf_64_clk _01052_ _00372_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_15847_ _01849_ _01850_ _01852_ _01858_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14558__A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11534__X _05423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18566_ clknet_leaf_13_clk _00986_ _00303_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[119\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13443__A1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15778_ game.CPU.applesa.ab.absxs.body_y\[105\] net446 vssd1 vssd1 vccd1 vccd1 _01790_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17517_ _02943_ _02944_ _02942_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11454__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14729_ _08559_ _08560_ net54 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__and3b_1
XFILLER_0_169_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18497_ net583 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__inv_2
XANTENNA__17185__A2 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19805__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17448_ net1258 _02772_ _02817_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__and3_1
XFILLER_0_184_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14564__Y game.CPU.walls.rand_wall.abduyd.next_wall\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19876__RESET_B net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18761__Q game.CPU.applesa.ab.absxs.body_x\[55\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ net1119 net1121 _02806_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__o21a_1
XANTENNA__13401__S net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12954__A0 _06757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19118_ net1182 _00158_ _00789_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[163\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09387__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19955__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12525__B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16696__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19049_ net1185 _00281_ _00720_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[94\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_357_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15836__B net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10045__B game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09834__B game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16999__A2 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14459__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout382_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_180_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09704_ net1150 game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1 vccd1
+ vccd1 _03947_ sky130_fd_sc_hd__xor2_1
XANTENNA__15852__A game.CPU.applesa.ab.absxs.body_y\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16300__X _02300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_241_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19335__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09850__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ net1148 game.CPU.applesa.ab.absxs.body_y\[17\] vssd1 vssd1 vccd1 vccd1 _03878_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout170_X net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1291_A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10996__A game.CPU.applesa.ab.absxs.body_y\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_222_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout647_A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09566_ net1144 game.CPU.applesa.ab.absxs.body_y\[77\] vssd1 vssd1 vccd1 vccd1 _03809_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_306_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19485__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout814_A game.CPU.applesa.ab.check_walls.above.walls\[70\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09497_ net1110 game.CPU.applesa.ab.check_walls.above.walls\[48\] vssd1 vssd1 vccd1
+ vccd1 _03740_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10799__A2 _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11996__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_322_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09996__S _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11996__B2 game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16923__A2 _02643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_322_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_286_Right_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_191_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18671__Q game.CPU.applesa.ab.absxs.body_y\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10410_ net1260 _04556_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__nand2_1
XANTENNA__09297__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11390_ _05275_ _05276_ _05277_ _05278_ _05264_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__a41o_1
XANTENNA__10507__Y _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16687__A1 _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10341_ _04338_ _04486_ _04508_ _04512_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__o211a_1
XFILLER_0_249_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14490__X _08364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18403__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13060_ game.writer.tracker.frame\[244\] game.writer.tracker.frame\[245\] net1027
+ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__mux2_1
X_10272_ net1171 _04367_ _04369_ game.CPU.applesa.ab.YMAX\[0\] vssd1 vssd1 vccd1 vccd1
+ _04465_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout971_X net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15746__B net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12722__Y _06596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12011_ game.CPU.applesa.ab.check_walls.above.walls\[76\] net554 vssd1 vssd1 vccd1
+ vccd1 _05898_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_280_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__B game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17100__A2 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13348__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_306_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09463__C net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13122__A0 game.writer.tracker.frame\[176\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19007__Q game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_245_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout460 net464 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_4
Xfanout471 net472 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_144_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15662__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16750_ net184 _02391_ net101 _02586_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[174\]
+ sky130_fd_sc_hd__a31o_1
Xfanout482 net486 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_4
Xfanout493 net494 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_4
X_13962_ net867 net784 _03478_ net960 _07835_ vssd1 vssd1 vccd1 vccd1 _07836_ sky130_fd_sc_hd__a221o_1
XANTENNA__09877__B1 _04118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16210__X _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15701_ game.CPU.applesa.ab.check_walls.above.walls\[156\] net342 vssd1 vssd1 vccd1
+ vccd1 _01713_ sky130_fd_sc_hd__or2_1
X_12913_ net509 _06786_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__or2_1
X_16681_ _02238_ _02555_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__nand2_8
XFILLER_0_220_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18702__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ net875 game.CPU.applesa.ab.check_walls.above.walls\[59\] _03415_ net952 vssd1
+ vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__19828__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18420_ net627 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__inv_2
X_15632_ _01636_ _01637_ _01638_ _01639_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__or4_1
X_12844_ _06714_ _06715_ _06717_ _06716_ net490 net682 vssd1 vssd1 vccd1 vccd1 _06718_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12228__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12859__S0 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14097__B net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18351_ net592 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ net576 _01581_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12775_ game.writer.tracker.frame\[128\] game.writer.tracker.frame\[129\] net1033
+ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_291_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17167__A2 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ net2019 net722 _02757_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[555\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_185_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14514_ _03207_ net1069 net861 game.CPU.apple_location2\[5\] _08384_ vssd1 vssd1
+ vccd1 vccd1 _08388_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11726_ net812 net301 _05611_ _05613_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__o211a_1
X_18282_ net622 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
X_15494_ _08040_ _08369_ _01471_ _01517_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__o31a_1
XANTENNA__18852__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17233_ _02418_ net123 net121 _02739_ net1575 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[504\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_232_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_253_Right_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14445_ _03263_ net1060 net861 game.CPU.applesa.ab.absxs.body_y\[89\] _08318_ vssd1
+ vssd1 vccd1 vccd1 _08319_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_330_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11657_ net829 net261 vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__nand2_1
X_17164_ _02456_ _02720_ net727 vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10608_ game.CPU.applesa.ab.absxs.body_x\[83\] _04673_ _04674_ game.CPU.applesa.ab.absxs.body_x\[79\]
+ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__a22o_1
XANTENNA__16127__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14376_ game.CPU.applesa.ab.absxs.body_x\[82\] net1053 vssd1 vssd1 vccd1 vccd1 _08250_
+ sky130_fd_sc_hd__xnor2_1
X_11588_ net564 _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__nor2_1
XANTENNA__09801__B1 game.CPU.applesa.ab.check_walls.above.walls\[106\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19208__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12345__B net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16115_ game.CPU.applesa.ab.absxs.body_x\[68\] net355 vssd1 vssd1 vccd1 vccd1 _02127_
+ sky130_fd_sc_hd__xnor2_1
X_13327_ _06725_ _06727_ _06734_ _06726_ net695 net476 vssd1 vssd1 vccd1 vccd1 _07201_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17095_ _02489_ net60 _02700_ net1651 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[405\]
+ sky130_fd_sc_hd__a22o_1
X_10539_ _03197_ _04606_ net850 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__a21o_2
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18313__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__A2_N net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09494__X _03737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16046_ _02050_ _02051_ _02053_ _02054_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__a22o_1
X_13258_ game.writer.tracker.frame\[454\] game.writer.tracker.frame\[455\] net1015
+ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__mux2_1
XANTENNA__15656__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_268_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12209_ game.CPU.applesa.ab.check_walls.above.walls\[143\] net422 vssd1 vssd1 vccd1
+ vccd1 _06095_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_244_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12361__A game.CPU.applesa.ab.absxs.body_x\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13189_ game.writer.tracker.frame\[434\] game.writer.tracker.frame\[435\] net1035
+ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__mux2_1
XANTENNA__19358__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11911__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19805_ clknet_leaf_38_clk game.writer.tracker.next_frame\[400\] net1328 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[400\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11911__B2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17997_ net637 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_166_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_257_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13113__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13744__X _07618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15672__A game.CPU.applesa.ab.check_walls.above.walls\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_19736_ clknet_leaf_15_clk game.writer.tracker.next_frame\[331\] net1289 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[331\] sky130_fd_sc_hd__dfrtp_1
X_16948_ _02394_ net86 net713 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__o21a_1
XFILLER_0_223_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16487__B _02434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13904__B net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10478__B2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18756__Q game.CPU.applesa.ab.absxs.body_x\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16879_ game.writer.tracker.frame\[258\] _02631_ vssd1 vssd1 vccd1 vccd1 _02632_
+ sky130_fd_sc_hd__and2_1
X_19667_ clknet_leaf_29_clk game.writer.tracker.next_frame\[262\] net1291 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[262\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16602__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16602__B2 game.writer.tracker.frame\[98\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09420_ net1098 _03261_ _03262_ net1107 _03657_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__a221o_1
X_18618_ clknet_leaf_13_clk _01035_ _00355_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[112\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_149_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19598_ clknet_leaf_35_clk game.writer.tracker.next_frame\[193\] net1346 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[193\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13416__A1 _07032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09351_ net1111 game.CPU.applesa.ab.absxs.body_x\[8\] vssd1 vssd1 vccd1 vccd1 _03594_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_47_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18549_ net615 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_255_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13920__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09282_ game.CPU.applesa.good_collision2 game.CPU.applesa.ab.good_collision vssd1
+ vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__or2_4
XFILLER_0_306_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_177_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_220_Right_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout130_A _02276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout228_A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13131__S net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11440__A game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14392__A2 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12255__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16669__B2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12970__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_344_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload70 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_fanout1137_A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout597_A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_266_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09564__B net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10705__A2 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17094__A1 _02237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20034__1382 vssd1 vssd1 vccd1 vccd1 net1382 _20034__1382/LO sky130_fd_sc_hd__conb_1
XFILLER_0_100_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09571__A2 game.CPU.applesa.ab.absxs.body_x\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16678__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ game.CPU.applesa.ab.absxs.body_x\[36\] vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__inv_2
XANTENNA__16841__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_355_Right_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout931_A _03190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19204__D _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_355_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09618_ net1150 game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 _03861_ sky130_fd_sc_hd__xor2_1
X_10890_ _04778_ _04790_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__xor2_1
XANTENNA__18875__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_333_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11334__B net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_277_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09549_ net1142 _03322_ game.CPU.applesa.ab.absxs.body_y\[113\] net899 _03791_ vssd1
+ vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__a221o_1
XANTENNA__14485__X _08359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19727__RESET_B net1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ _06432_ _06433_ _06434_ _06436_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__or4_1
XFILLER_0_65_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10641__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11511_ game.CPU.applesa.ab.check_walls.above.walls\[1\] net772 vssd1 vssd1 vccd1
+ vccd1 _05400_ sky130_fd_sc_hd__xor2_1
XANTENNA__09739__B game.CPU.applesa.ab.check_walls.above.walls\[65\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12491_ game.CPU.applesa.ab.absxs.body_y\[80\] net359 vssd1 vssd1 vccd1 vccd1 _06368_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11548__A1_N net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14230_ _08098_ _08099_ _08102_ _08103_ vssd1 vssd1 vccd1 vccd1 _08104_ sky130_fd_sc_hd__a22o_1
XANTENNA__14383__A2 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11442_ net825 net261 _05328_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13040__C1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_297_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12165__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14161_ net1094 net879 net874 net1087 _08034_ vssd1 vssd1 vccd1 vccd1 _08035_ sky130_fd_sc_hd__a221o_1
X_11373_ game.CPU.applesa.ab.check_walls.above.walls\[38\] net256 _05256_ net565 _05261_
+ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__a221o_1
XFILLER_0_296_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16205__X _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13112_ game.writer.tracker.frame\[140\] game.writer.tracker.frame\[141\] net991
+ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__mux2_1
X_10324_ net1933 _04500_ vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_308_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19500__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09755__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14092_ net961 net830 vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__xor2_1
XFILLER_0_277_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17609__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13043_ _06872_ _06887_ net697 vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__mux2_1
XANTENNA__14540__C1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10255_ net759 net571 _04447_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a21oi_1
X_17920_ net604 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__inv_2
XFILLER_0_265_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13894__A1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1200 net1201 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__buf_1
XANTENNA__13894__B2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17085__A1 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1211 net1212 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_2
X_17851_ game.writer.updater.commands.count\[10\] _03169_ _03175_ vssd1 vssd1 vccd1
+ vccd1 _03176_ sky130_fd_sc_hd__o21ai_1
X_10186_ _04368_ _04373_ _04376_ _04378_ _04377_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__a221o_1
Xfanout1222 net1224 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__clkbuf_2
Xfanout1233 net1234 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__clkbuf_2
Xfanout1244 net1246 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__clkbuf_2
XANTENNA__19650__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16802_ _02487_ net104 _02601_ net1845 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[211\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16832__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1255 net1256 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__clkbuf_2
X_17782_ game.CPU.applesa.twoapples.count\[1\] game.CPU.applesa.twoapples.count\[0\]
+ net1163 game.CPU.applesa.twoapples.count\[2\] vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__a31o_1
Xfanout1266 game.CPU.applesa.ab.absxs.body_x\[101\] vssd1 vssd1 vccd1 vccd1 net1266
+ sky130_fd_sc_hd__buf_4
XFILLER_0_205_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14994_ net1223 net1251 game.CPU.applesa.ab.check_walls.above.walls\[22\] vssd1 vssd1
+ vccd1 vccd1 _00211_ sky130_fd_sc_hd__and3_1
Xfanout1277 net1278 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__clkbuf_2
Xfanout1288 net1290 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__clkbuf_4
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_4
Xfanout1299 net1300 vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__clkbuf_4
X_19521_ clknet_leaf_21_clk game.writer.tracker.next_frame\[116\] net1335 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[116\] sky130_fd_sc_hd__dfrtp_1
X_16733_ _02364_ net101 _02580_ net1699 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[163\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18576__Q game.CPU.applesa.ab.absxs.body_y\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13945_ net875 game.CPU.applesa.ab.check_walls.above.walls\[67\] _03419_ net965 _07814_
+ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__a221o_1
XFILLER_0_205_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14413__A1_N game.CPU.applesa.ab.absxs.body_x\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_322_Right_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_64_clk_X clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19452_ clknet_leaf_47_clk game.writer.tracker.next_frame\[47\] net1295 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[47\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload6_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16664_ net2040 _02548_ _02549_ net128 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[125\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_319_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13876_ _07746_ _07747_ _07748_ _07749_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__and4_1
XFILLER_0_201_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_243_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18403_ net618 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__inv_2
X_15615_ game.CPU.applesa.ab.check_walls.above.walls\[82\] net469 vssd1 vssd1 vccd1
+ vccd1 _01627_ sky130_fd_sc_hd__xnor2_1
X_12827_ net176 vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__inv_2
XANTENNA__11244__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19383_ clknet_leaf_3_clk _01389_ _00963_ vssd1 vssd1 vccd1 vccd1 game.CPU.bodymain1.main.score\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_16595_ net113 _02509_ net716 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__o21a_1
XFILLER_0_347_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18334_ net599 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15546_ _01565_ _01566_ _01557_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__a21o_1
XFILLER_0_173_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12758_ _06579_ _06585_ _06584_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16899__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11709_ _05473_ _05534_ _05566_ _05597_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__and4_1
X_18265_ net645 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
XANTENNA__11290__D1 _05084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15477_ _01459_ _01484_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12689_ net1065 net1057 _06550_ _06562_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__o22a_2
XFILLER_0_71_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12356__A game.CPU.applesa.ab.absxs.body_x\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17216_ _02238_ _02241_ _02520_ _02619_ net713 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__o41a_1
XFILLER_0_115_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ game.CPU.applesa.ab.absxs.body_x\[26\] net880 net857 game.CPU.applesa.ab.absxs.body_y\[27\]
+ vssd1 vssd1 vccd1 vccd1 _08302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_343_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18196_ net581 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_250_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17147_ _02422_ net58 _02716_ net1716 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[441\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14359_ game.CPU.applesa.ab.absxs.body_y\[102\] net951 vssd1 vssd1 vccd1 vccd1 _08233_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__14571__A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17312__A2 _02535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_268_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19180__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09665__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17078_ _02291_ _02693_ net735 vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18748__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12137__A1 game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_338_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12137__B2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16029_ game.CPU.applesa.ab.absxs.body_y\[95\] net432 net445 game.CPU.applesa.ab.absxs.body_y\[93\]
+ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__15874__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10163__X _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17076__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10699__A1 game.CPU.applesa.ab.absxs.body_y\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10699__B2 game.CPU.applesa.ab.absxs.body_y\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_236_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13915__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19719_ clknet_leaf_35_clk game.writer.tracker.next_frame\[314\] net1345 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[314\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11962__A2_N net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16010__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11435__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16587__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09403_ net922 game.CPU.applesa.ab.check_walls.above.walls\[90\] net807 net895 _03640_
+ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__o221a_1
XANTENNA__12965__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_A game.CPU.walls.rand_wall.abduyd.next_wall\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _03571_ _03576_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__or2_1
XANTENNA__12612__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14465__B net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10993__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17000__A1 _02322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_319_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11820__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ game.CPU.randy.counter1.count1\[3\] vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_350_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout512_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1254_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11170__A net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_279_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19523__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09196_ game.CPU.applesa.ab.check_walls.above.walls\[122\] vssd1 vssd1 vccd1 vccd1
+ _03445_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16680__B net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_279_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_214_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1042_X net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout881_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_248_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout979_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19673__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17792__A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1307_X net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10040_ net1171 _04218_ _04220_ game.CPU.applesa.ab.YMAX\[0\] vssd1 vssd1 vccd1 vccd1
+ _04248_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11329__B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19780__Q game.writer.tracker.frame\[375\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 game.CPU.up_button.eD1.D vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 game.CPU.walls.abc.number\[3\] vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold32 game.CPU.applesa.twomode.number\[3\] vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_303_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold43 game.CPU.applesa.twomode.number\[2\] vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold54 game.CPU.randy.f1.a1.count\[13\] vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_279_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold65 game.CPU.applesa.ab.apple_location\[1\] vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 net45 vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 game.writer.tracker.frame\[330\] vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold98 game.writer.tracker.frame\[263\] vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11991_ _05319_ _05323_ _05877_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__or3_1
X_13730_ game.writer.tracker.frame\[223\] net710 net673 game.writer.tracker.frame\[224\]
+ vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__o22a_1
XFILLER_0_242_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10942_ game.CPU.applesa.ab.absxs.body_y\[29\] net405 vssd1 vssd1 vccd1 vccd1 _04832_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_344_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_356_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11064__B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19053__CLK net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13661_ game.writer.tracker.frame\[13\] game.writer.tracker.frame\[15\] game.writer.tracker.frame\[16\]
+ game.writer.tracker.frame\[14\] net971 net1004 vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__mux4_1
X_10873_ game.CPU.applesa.ab.apple_possible\[4\] net759 vssd1 vssd1 vccd1 vccd1 _04775_
+ sky130_fd_sc_hd__or2_2
XANTENNA__14053__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14053__B2 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15400_ game.writer.updater.commands.count\[11\] game.writer.updater.commands.count\[10\]
+ game.writer.updater.commands.count\[12\] vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__a21o_1
XANTENNA__13560__A net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12612_ game.CPU.applesa.ab.absxs.body_y\[21\] net523 net359 game.CPU.applesa.ab.absxs.body_y\[20\]
+ _06457_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__a221o_1
X_16380_ net172 _02357_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__nor2_1
XANTENNA__13800__A1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13592_ _07464_ _07465_ net509 vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_197_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10614__A1 game.CPU.applesa.ab.absxs.body_x\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15331_ game.CPU.applesa.twomode.number\[7\] _08870_ _00029_ vssd1 vssd1 vccd1 vccd1
+ _08874_ sky130_fd_sc_hd__a21oi_1
XANTENNA__17967__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12543_ game.CPU.applesa.ab.absxs.body_y\[43\] net367 vssd1 vssd1 vccd1 vccd1 _06420_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__09480__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10248__X _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19020__Q game.CPU.applesa.ab.check_walls.above.walls\[65\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_314_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09480__B2 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18050_ net661 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15262_ _08818_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__inv_2
XFILLER_0_325_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12474_ game.CPU.applesa.ab.absxs.body_y\[58\] net520 vssd1 vssd1 vccd1 vccd1 _06351_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_340_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17001_ _02486_ net83 _02672_ net2025 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[339\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_289_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14213_ game.CPU.applesa.ab.absxs.body_y\[95\] net939 vssd1 vssd1 vccd1 vccd1 _08087_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11425_ _05292_ _05295_ _05313_ _05279_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__a211o_1
X_15193_ _04586_ _08761_ _08762_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__a21o_1
XANTENNA_7 _02179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14144_ _07907_ _07908_ _07913_ _07915_ net358 vssd1 vssd1 vccd1 vccd1 _08018_ sky130_fd_sc_hd__a41o_1
XFILLER_0_284_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11356_ game.CPU.applesa.ab.check_walls.above.walls\[143\] net258 vssd1 vssd1 vccd1
+ vccd1 _05245_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_78_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13316__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15856__A2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ game.CPU.randy.f1.a1.count\[6\] game.CPU.randy.f1.a1.count\[5\] _04489_ vssd1
+ vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__and3_1
X_14075_ _07943_ _07946_ _07947_ _07948_ vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__and4_1
X_18952_ clknet_leaf_68_clk net1409 _00623_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13867__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11287_ _04982_ _04983_ _04989_ _04990_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a22o_1
XANTENNA__17058__A1 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13026_ _06862_ _06881_ net697 vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_253_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17903_ net669 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__inv_2
XANTENNA__11239__B net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10238_ _04392_ _04399_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__nand2_1
XANTENNA__15934__B net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18883_ clknet_leaf_7_clk game.CPU.randy.f1.c1.innerCount\[13\] _00578_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[13\] sky130_fd_sc_hd__dfrtp_1
Xfanout1030 net1034 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16805__A1 _02490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 net1042 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__buf_4
XFILLER_0_280_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17834_ game.writer.updater.commands.count\[6\] _03161_ vssd1 vssd1 vccd1 vccd1 _03163_
+ sky130_fd_sc_hd__nand2_1
Xfanout1052 net1053 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__clkbuf_4
X_10169_ net1168 game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1 vccd1 vccd1 _04362_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_163_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1063 net1068 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__buf_4
Xfanout1074 net1077 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__buf_4
XFILLER_0_89_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1085 net1087 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__buf_4
Xfanout1096 net1097 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_4
X_14977_ net1226 net1253 game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1
+ vccd1 vccd1 _00132_ sky130_fd_sc_hd__and3_1
X_17765_ _03109_ _03118_ _03119_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__and3_1
XANTENNA__19649__RESET_B net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19504_ clknet_leaf_29_clk game.writer.tracker.next_frame\[99\] net1283 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[99\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16716_ net1840 _02572_ _02573_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[153\]
+ sky130_fd_sc_hd__a21o_1
X_20010__1379 vssd1 vssd1 vccd1 vccd1 net1379 _20010__1379/LO sky130_fd_sc_hd__conb_1
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13928_ net1063 game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1 vssd1 vccd1
+ vccd1 _07802_ sky130_fd_sc_hd__nand2_1
X_17696_ game.CPU.walls.rand_wall.count\[0\] net1175 vssd1 vssd1 vccd1 vccd1 _03075_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_254_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_297_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17230__A1 _02415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16647_ net1810 _02540_ _02542_ net126 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[115\]
+ sky130_fd_sc_hd__a22o_1
X_19435_ clknet_leaf_41_clk game.writer.tracker.next_frame\[30\] net1332 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13859_ game.writer.tracker.frame\[554\] net842 net835 game.writer.tracker.frame\[553\]
+ net281 vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_44_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12638__X _06515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13470__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16578_ _02301_ _02493_ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_252_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19366_ clknet_leaf_68_clk _01372_ _00947_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_186_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15529_ net1065 net1049 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__xor2_1
X_18317_ net615 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__inv_2
XANTENNA__09379__B net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19297_ clknet_leaf_68_clk net323 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.x_final\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_20033__1381 vssd1 vssd1 vccd1 vccd1 net1381 _20033__1381/LO sky130_fd_sc_hd__conb_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09050_ game.CPU.applesa.ab.absxs.body_y\[79\] vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__inv_2
X_18248_ net644 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_59_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10620__A4 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18570__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19696__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18179_ net608 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__inv_2
Xhold502 game.writer.tracker.frame\[12\] vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_349_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold513 game.writer.tracker.frame\[570\] vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold524 game.writer.tracker.frame\[10\] vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09774__A2 game.CPU.applesa.ab.YMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 game.writer.tracker.frame\[69\] vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 game.CPU.walls.rand_wall.count_luck\[6\] vssd1 vssd1 vccd1 vccd1 net1931
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 game.writer.tracker.frame\[189\] vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16005__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold568 game.writer.tracker.frame\[158\] vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold579 game.writer.tracker.frame\[521\] vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ net1122 _04172_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__or2_1
XANTENNA__10334__A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_263_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17049__A1 _02415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11149__B net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ _03674_ _03675_ _03916_ _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__o211a_1
XANTENNA__15844__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_A _05858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12530__A1 game.CPU.applesa.ab.absxs.body_x\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10988__B game.CPU.applesa.ab.absxs.next_head\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19076__CLK net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19105__Q game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout462_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_352_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17221__A1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_338_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout250_X net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout727_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16575__A3 _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_274_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_314_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16980__B1 _02665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_216_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09317_ net1140 game.CPU.applesa.ab.absxs.body_y\[66\] vssd1 vssd1 vccd1 vccd1 _03560_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11612__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18913__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1257_X net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14338__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ game.CPU.randy.counter1.count1\[17\] vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__inv_2
XFILLER_0_334_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_330_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09179_ game.CPU.applesa.ab.check_walls.above.walls\[89\] vssd1 vssd1 vccd1 vccd1
+ _03428_ sky130_fd_sc_hd__inv_2
XANTENNA__13641__S0 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12724__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17288__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ game.CPU.applesa.ab.absxs.body_x\[95\] net408 vssd1 vssd1 vccd1 vccd1 _05100_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12190_ game.CPU.applesa.ab.check_walls.above.walls\[126\] net417 vssd1 vssd1 vccd1
+ vccd1 _06076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_266_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout884_X net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput11 net11 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_0_31_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput9 net9 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XANTENNA__11854__A2_N net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
X_11141_ _05020_ _05029_ _05030_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_285_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_227_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11072_ _04954_ _04959_ _04960_ _04961_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__or4_2
XFILLER_0_290_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15754__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14510__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19419__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ _04230_ _04229_ _04227_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__or3b_1
X_14900_ _08673_ _08676_ vssd1 vssd1 vccd1 vccd1 _08677_ sky130_fd_sc_hd__and2_1
XANTENNA__09752__B net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15880_ net791 net438 vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__nor2_1
XANTENNA__10531__X _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14831_ _08632_ vssd1 vssd1 vccd1 vccd1 _08633_ sky130_fd_sc_hd__inv_2
XANTENNA__14274__A1 game.CPU.applesa.ab.absxs.body_x\[49\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_355_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_291_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14274__B2 game.CPU.applesa.ab.absxs.body_x\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11075__A game.CPU.applesa.ab.absxs.body_x\[40\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15770__A game.CPU.applesa.ab.absxs.body_y\[106\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_203_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17550_ net1271 _02778_ net428 _02973_ _02975_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_199_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ game.CPU.randy.counter1.count\[11\] net265 vssd1 vssd1 vccd1 vccd1 _08583_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__19569__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ _05193_ _05860_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__and2_1
X_16501_ _02345_ _02445_ net730 vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__o21a_1
X_13713_ game.writer.tracker.frame\[201\] game.writer.tracker.frame\[203\] game.writer.tracker.frame\[204\]
+ game.writer.tracker.frame\[202\] net974 net1011 vssd1 vssd1 vccd1 vccd1 _07587_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_316_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _04375_ _04472_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__or2_1
X_17481_ _02901_ _02909_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_224_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14026__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14693_ game.CPU.randy.counter1.count1\[12\] _08530_ _08529_ vssd1 vssd1 vccd1 vccd1
+ _08532_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14026__B2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16432_ net134 net114 _02394_ net724 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__o31a_1
XFILLER_0_195_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19220_ clknet_leaf_69_clk _01314_ _00859_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_location\[2\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11803__A game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13644_ game.writer.tracker.frame\[30\] net845 net838 game.writer.tracker.frame\[29\]
+ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__o22a_1
XFILLER_0_224_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10856_ _03500_ game.CPU.randy.counter1.count1\[13\] game.CPU.randy.counter1.count1\[12\]
+ _03501_ _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a221o_1
XFILLER_0_160_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18593__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19151_ net1187 _00194_ _00822_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[196\]
+ sky130_fd_sc_hd__dfrtp_4
X_16363_ net1984 net737 _02346_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[27\]
+ sky130_fd_sc_hd__and3_1
X_13575_ game.writer.tracker.frame\[321\] game.writer.tracker.frame\[323\] game.writer.tracker.frame\[324\]
+ game.writer.tracker.frame\[322\] net979 net1030 vssd1 vssd1 vccd1 vccd1 _07449_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10787_ game.CPU.applesa.ab.absxs.body_y\[50\] _04630_ vssd1 vssd1 vccd1 vccd1 _04725_
+ sky130_fd_sc_hd__and2_1
X_18102_ net603 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__inv_2
XFILLER_0_240_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15314_ game.CPU.applesa.twomode.number\[4\] _08854_ vssd1 vssd1 vccd1 vccd1 _08860_
+ sky130_fd_sc_hd__nand2_1
X_19082_ net1185 _00118_ _00753_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[127\]
+ sky130_fd_sc_hd__dfrtp_4
X_12526_ game.CPU.applesa.ab.absxs.body_x\[96\] net381 vssd1 vssd1 vccd1 vccd1 _06403_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16294_ net1008 _08400_ _02261_ net971 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15929__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13537__A0 game.writer.tracker.frame\[81\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_240_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18033_ net601 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
X_15245_ game.CPU.kyle.L1.cnt_500hz\[6\] game.CPU.kyle.L1.cnt_500hz\[9\] vssd1 vssd1
+ vccd1 vccd1 _08806_ sky130_fd_sc_hd__nor2_1
X_12457_ net1269 net377 net360 game.CPU.applesa.ab.absxs.body_y\[48\] _06333_ vssd1
+ vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__o221a_1
XFILLER_0_340_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17279__A1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15010__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ net799 net251 vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__nand2_1
X_15176_ game.CPU.bodymain1.main.score\[7\] net1115 net1114 vssd1 vssd1 vccd1 vccd1
+ _08752_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_327_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12388_ _03348_ game.CPU.applesa.twoapples.absxs.next_head\[7\] vssd1 vssd1 vccd1
+ vccd1 _06265_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12353__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__A1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14127_ net1075 _03390_ game.CPU.applesa.ab.check_walls.above.walls\[27\] net875
+ _07998_ vssd1 vssd1 vccd1 vccd1 _08001_ sky130_fd_sc_hd__o221a_1
X_11339_ net775 _05227_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12921__X _06795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19984_ clknet_leaf_46_clk _01408_ net1280 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.y\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_18935_ clknet_leaf_14_clk net1404 net1282 vssd1 vssd1 vccd1 vccd1 game.CPU.reset_button1.eD1.Q2
+ sky130_fd_sc_hd__dfrtp_1
X_14058_ net958 game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1 vccd1
+ vccd1 _07932_ sky130_fd_sc_hd__xor2_1
XFILLER_0_281_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12512__A1 game.CPU.applesa.ab.absxs.body_y\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13009_ game.writer.tracker.frame\[552\] game.writer.tracker.frame\[553\] net1006
+ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_253_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12512__B2 game.CPU.applesa.ab.absxs.body_y\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18866_ clknet_leaf_0_clk _01257_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_17817_ game.writer.updater.commands.count\[1\] game.writer.updater.commands.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__nand2_1
XFILLER_0_265_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18797_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[0\] _00534_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14265__B2 game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_206_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15680__A game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17748_ _04255_ _04252_ net1162 vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_338_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14567__Y game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17203__A1 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18936__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14296__A game.CPU.applesa.ab.absxs.body_x\[53\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17679_ _03062_ _03065_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13404__S net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15603__A1_N game.CPU.applesa.ab.check_walls.above.walls\[113\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19418_ clknet_leaf_48_clk game.writer.tracker.next_frame\[13\] net1303 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_336_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_335_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11432__B net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19349_ clknet_leaf_70_clk net369 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.y_final\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_351_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09102_ game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__inv_2
XANTENNA__17400__A _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11251__B2 game.CPU.applesa.ab.absxs.body_x\[115\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16714__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_304_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_198_Right_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15839__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10048__B net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13199__X _07073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_288_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09033_ game.CPU.applesa.ab.absxs.body_x\[19\] vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__inv_2
XFILLER_0_331_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout210_A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13623__S0 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout308_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_211_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold310 game.writer.tracker.frame\[503\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_248_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold321 game.writer.tracker.frame\[52\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_300_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold332 game.writer.tracker.frame\[266\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12263__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold343 game.writer.tracker.frame\[301\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold354 game.writer.tracker.frame\[213\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold365 game.CPU.applesa.steady\[0\] vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 game.writer.tracker.frame\[379\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10762__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 game.writer.tracker.frame\[445\] vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_6_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1217_A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold398 game.writer.tracker.frame\[315\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 game.CPU.applesa.ab.check_walls.above.walls\[110\] vssd1 vssd1 vccd1 vccd1
+ net801 sky130_fd_sc_hd__buf_2
XFILLER_0_284_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09935_ net1121 net1124 vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__and2_1
Xfanout812 game.CPU.applesa.ab.check_walls.above.walls\[78\] vssd1 vssd1 vccd1 vccd1
+ net812 sky130_fd_sc_hd__clkbuf_4
Xfanout823 game.CPU.applesa.ab.check_walls.above.walls\[37\] vssd1 vssd1 vccd1 vccd1
+ net823 sky130_fd_sc_hd__clkbuf_4
Xfanout834 net840 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__buf_4
XANTENNA__10999__A game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_272_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout677_A _06600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 _06574_ vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_4
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20055_ net1373 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_256_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout856 net857 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_4
X_09866_ net1142 game.CPU.applesa.ab.absxs.body_y\[110\] vssd1 vssd1 vccd1 vccd1 _04109_
+ sky130_fd_sc_hd__xor2_1
Xfanout867 net868 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1005_X net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10514__B1 _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout878 net879 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_13_Left_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19711__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout889 _03368_ vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09380__B1 _03385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_300_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12599__A2_N net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout844_A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ net922 game.CPU.applesa.ab.absxs.body_x\[42\] game.CPU.applesa.ab.absxs.body_y\[40\]
+ net895 _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14256__B2 game.CPU.applesa.ab.absxs.body_x\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17134__X _02713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_222_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09999__S _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18674__Q game.CPU.applesa.ab.absxs.body_x\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14008__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09683__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14008__B2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19861__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10710_ game.CPU.applesa.ab.absxs.body_y\[62\] net425 _04711_ net934 vssd1 vssd1
+ vccd1 vccd1 _01069_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_339_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11690_ net817 net252 vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13767__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_341_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10641_ net932 game.CPU.applesa.ab.absxs.body_x\[44\] net561 _04688_ vssd1 vssd1
+ vccd1 vccd1 _01115_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_194_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Left_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_341_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13360_ _07230_ _07233_ net229 vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_311_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10572_ _03252_ net234 vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__nor2_1
XANTENNA__15749__B net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_307_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12311_ game.CPU.applesa.ab.check_walls.above.walls\[191\] net421 vssd1 vssd1 vccd1
+ vccd1 _06197_ sky130_fd_sc_hd__nand2_1
X_13291_ _06763_ _06764_ _06779_ _06765_ net705 net497 vssd1 vssd1 vccd1 vccd1 _07165_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09747__B game.CPU.applesa.ab.check_walls.above.walls\[68\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15030_ net1222 net1256 game.CPU.applesa.ab.check_walls.above.walls\[58\] vssd1 vssd1
+ vccd1 vccd1 _00250_ sky130_fd_sc_hd__and3_1
XFILLER_0_310_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12242_ _06124_ _06127_ _06125_ _06126_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__or4b_1
XANTENNA__14192__B1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12173__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12173_ net807 net554 vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17130__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16213__X _02225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19994__RESET_B net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09763__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124_ game.CPU.applesa.ab.absxs.body_y\[16\] net534 vssd1 vssd1 vccd1 vccd1 _05014_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_263_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16981_ net190 _02460_ net91 _02665_ net1519 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[326\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_275_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19923__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Left_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18720_ clknet_leaf_69_clk _01137_ _00457_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[90\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17980__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11055_ game.CPU.applesa.ab.absxs.body_y\[105\] net542 net539 game.CPU.applesa.ab.absxs.body_y\[106\]
+ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a2bb2o_1
X_15932_ game.CPU.applesa.ab.check_walls.above.walls\[120\] net354 vssd1 vssd1 vccd1
+ vccd1 _01944_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_147_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_322_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20032__1380 vssd1 vssd1 vccd1 vccd1 net1380 _20032__1380/LO sky130_fd_sc_hd__conb_1
XANTENNA__19391__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ net910 _04212_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__xnor2_2
X_18651_ clknet_leaf_51_clk _01068_ _00388_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[61\]
+ sky130_fd_sc_hd__dfrtp_4
X_15863_ game.CPU.applesa.ab.absxs.body_x\[114\] net467 vssd1 vssd1 vccd1 vccd1 _01875_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__18959__CLK net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__B _04563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14814_ game.CPU.randy.counter1.count\[13\] _08621_ net138 vssd1 vssd1 vccd1 vccd1
+ _08623_ sky130_fd_sc_hd__o21ai_1
X_17602_ _03009_ _03017_ net582 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_349_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13455__C1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18582_ clknet_leaf_53_clk _01002_ _00319_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[43\]
+ sky130_fd_sc_hd__dfrtp_4
X_15794_ game.CPU.applesa.ab.absxs.body_x\[48\] net355 net433 game.CPU.applesa.ab.absxs.body_y\[51\]
+ _01805_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__o221a_1
XFILLER_0_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10808__A1 game.CPU.applesa.ab.absxs.body_y\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17533_ net1119 _02939_ _02945_ _02960_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__a211o_1
X_14745_ game.CPU.randy.counter1.count1\[14\] game.CPU.randy.counter1.count1\[13\]
+ _08567_ vssd1 vssd1 vccd1 vccd1 _08571_ sky130_fd_sc_hd__and3_1
X_11957_ net815 net309 net303 net814 vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__a22oi_1
XANTENNA__17540__A_N _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_294_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10908_ net1243 game.CPU.applesa.enable_in _04734_ vssd1 vssd1 vccd1 vccd1 _00010_
+ sky130_fd_sc_hd__mux2_1
X_17464_ _02886_ _02892_ _02890_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__o21a_1
XANTENNA__11481__A1 _04450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15005__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14676_ game.CPU.randy.counter1.count1\[3\] _04356_ vssd1 vssd1 vccd1 vccd1 _08515_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_317_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11888_ net751 _05350_ net394 game.CPU.applesa.ab.check_walls.above.walls\[20\] _05774_
+ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__o221a_1
XANTENNA__12348__B net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13758__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16415_ net1683 _02380_ _02383_ net135 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[42\]
+ sky130_fd_sc_hd__a22o_1
X_19203_ clknet_leaf_70_clk _00016_ _00851_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.XMAX\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_345_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13627_ _07499_ _07500_ net514 vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10839_ _03511_ game.CPU.randy.counter1.count\[4\] _03509_ game.CPU.randy.counter1.count1\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__a2bb2o_1
X_17395_ _03218_ game.CPU.kyle.L1.nextState\[0\] vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__nor2_4
XFILLER_0_116_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16346_ _06572_ _06573_ _06607_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__and3_1
X_19134_ net1184 _00175_ _00805_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[179\]
+ sky130_fd_sc_hd__dfrtp_4
X_13558_ game.writer.tracker.frame\[99\] net709 net834 game.writer.tracker.frame\[97\]
+ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__o22a_1
XANTENNA__12430__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15659__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12981__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19065_ net1190 _00100_ _00736_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_12509_ game.CPU.applesa.ab.absxs.body_x\[73\] net377 vssd1 vssd1 vccd1 vccd1 _06386_
+ sky130_fd_sc_hd__xnor2_1
X_16277_ net2047 net718 _02281_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[6\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_11_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16172__A1 game.CPU.applesa.ab.absxs.body_x\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13489_ _07117_ _07118_ _07144_ _07119_ net700 net487 vssd1 vssd1 vccd1 vccd1 _07363_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15228_ _08792_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14183__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18016_ net640 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__inv_2
XFILLER_0_298_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12083__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15675__A game.CPU.applesa.ab.check_walls.above.walls\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15159_ net1213 net1240 game.CPU.applesa.ab.check_walls.above.walls\[187\] vssd1
+ vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__and3_1
XANTENNA__17121__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_247_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16475__A2 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout108 net109 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_4
XANTENNA__19734__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_238_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18759__Q game.CPU.applesa.ab.absxs.body_x\[53\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19967_ clknet_leaf_41_clk game.writer.tracker.next_frame\[562\] net1326 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[562\] sky130_fd_sc_hd__dfrtp_1
Xfanout119 net120 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13907__B game.CPU.applesa.ab.check_walls.above.walls\[123\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_254_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09720_ net1106 game.CPU.applesa.ab.absxs.body_x\[84\] vssd1 vssd1 vccd1 vccd1 _03963_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__17890__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18918_ clknet_leaf_5_clk net1387 _00602_ vssd1 vssd1 vccd1 vccd1 game.CPU.down_button.eD1.Q1
+ sky130_fd_sc_hd__dfrtp_1
X_19898_ clknet_leaf_15_clk game.writer.tracker.next_frame\[493\] net1288 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[493\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09898__D1 _03577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ net1154 net785 vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__or2_1
XANTENNA__11427__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18849_ clknet_leaf_6_clk _01240_ _00559_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_124_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19884__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09582_ _03816_ _03820_ _03823_ _03824_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__or4_2
XANTENNA__13446__C1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_267_Right_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17114__B net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17188__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _05195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11443__A game.CPU.applesa.ab.check_walls.above.walls\[74\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_258_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11472__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16935__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_271_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12258__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11162__B game.CPU.applesa.ab.absxs.next_head\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12973__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12826__X _06700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout425_A _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_308_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1167_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16950__A3 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12421__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12972__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19264__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1334_A net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14174__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09016_ game.CPU.applesa.ab.absxs.body_x\[82\] vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_347_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold140 game.writer.tracker.frame\[233\] vssd1 vssd1 vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 game.writer.tracker.frame\[150\] vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_269_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12561__X _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold162 game.writer.tracker.frame\[143\] vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__B1 _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold173 game.writer.tracker.frame\[384\] vssd1 vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09583__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16466__A2 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_282_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold184 game.writer.tracker.frame\[515\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 game.writer.tracker.frame\[413\] vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout961_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_256_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12721__B _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 net623 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_224_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14477__B2 game.CPU.applesa.ab.absxs.body_y\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout631 net632 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_4
X_09918_ net1084 _04155_ _04159_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__a21oi_1
Xfanout642 net646 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_298_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout653 net655 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_2
XANTENNA_fanout73_A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout664 net667 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_4
Xfanout675 _07401_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14121__A1_N net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09353__B1 game.CPU.applesa.ab.absxs.body_y\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout686 net691 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_4
X_20038_ net1362 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
Xfanout697 net699 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_4
X_09849_ net1096 _03248_ _03314_ net1126 _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__a221o_1
XANTENNA__11337__B net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14488__X _08362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16847__C net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_358_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ game.writer.tracker.frame\[264\] game.writer.tracker.frame\[265\] net996
+ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_358_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_234_Right_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11811_ _05690_ _05696_ _05698_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_17_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ game.writer.tracker.frame\[378\] game.writer.tracker.frame\[379\] net1032
+ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09656__A1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13452__A2 _07321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09656__B2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13044__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14530_ _08028_ _08039_ vssd1 vssd1 vccd1 vccd1 _08404_ sky130_fd_sc_hd__or2_2
X_11742_ net572 _05523_ _05528_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_352_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14461_ _08325_ _08329_ _08330_ _08334_ vssd1 vssd1 vccd1 vccd1 _08335_ sky130_fd_sc_hd__or4_1
XANTENNA__19607__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11673_ net795 net314 vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__nand2_1
XFILLER_0_315_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12736__X _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16200_ _03270_ net344 net441 game.CPU.applesa.ab.absxs.body_y\[58\] _02211_ vssd1
+ vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__a221o_1
X_13412_ net484 _07283_ _07285_ net225 vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__a211o_1
X_17180_ net174 net144 _02479_ _02634_ net728 vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__o41a_1
X_10624_ game.CPU.applesa.ab.absxs.body_x\[65\] _04679_ _04680_ game.CPU.applesa.ab.absxs.body_x\[61\]
+ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__a22o_1
XANTENNA__09758__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12412__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14392_ _03223_ net1046 net863 game.CPU.applesa.ab.absxs.body_y\[5\] _08261_ vssd1
+ vssd1 vccd1 vccd1 _08266_ sky130_fd_sc_hd__a221o_1
X_16131_ _01753_ _01754_ _01755_ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__or4_1
XANTENNA__11766__A2 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13343_ net201 _07216_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__or2_1
X_10555_ _03281_ net330 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__nor2_1
XANTENNA__12184__A game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19757__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16062_ _03484_ net353 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__xnor2_1
XANTENNA__18631__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13274_ game.writer.tracker.frame\[494\] game.writer.tracker.frame\[495\] net997
+ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_267_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ game.CPU.applesa.ab.absxs.body_x\[86\] _04610_ _04611_ game.CPU.applesa.ab.absxs.body_x\[82\]
+ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__a22o_1
XFILLER_0_322_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15013_ net1220 net1249 game.CPU.applesa.ab.check_walls.above.walls\[41\] vssd1 vssd1
+ vccd1 vccd1 _00231_ sky130_fd_sc_hd__and3_1
XANTENNA__15495__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12225_ _05897_ _05898_ _06109_ _06110_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_324_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19821_ clknet_leaf_37_clk game.writer.tracker.next_frame\[416\] net1350 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[416\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_208_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12156_ net824 net553 vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16103__B net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ game.CPU.applesa.ab.absxs.body_x\[32\] net326 vssd1 vssd1 vccd1 vccd1 _04997_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__10741__A3 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19752_ clknet_leaf_25_clk game.writer.tracker.next_frame\[347\] net1322 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[347\] sky130_fd_sc_hd__dfrtp_1
X_16964_ _02425_ _02636_ net729 vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__o21a_1
X_12087_ net827 net297 vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__or2_1
XANTENNA__13140__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_271_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18703_ clknet_leaf_31_clk _01120_ _00440_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[57\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_88_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11038_ _04922_ _04925_ _04926_ _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__or4_1
X_15915_ net792 net336 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__nand2_1
XANTENNA__11247__B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19683_ clknet_leaf_35_clk game.writer.tracker.next_frame\[278\] net1338 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[278\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15942__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16895_ _02466_ net93 _02640_ net1758 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[265\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11151__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13691__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18634_ clknet_leaf_61_clk _01051_ _00371_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15846_ _01851_ _01853_ _01855_ _01857_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__or4_1
XFILLER_0_91_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11055__A2_N net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_201_Right_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18565_ clknet_leaf_13_clk _00985_ _00302_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[118\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_176_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09647__A1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_335_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ game.writer.tracker.frame\[558\] game.writer.tracker.frame\[559\] net1007
+ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__mux2_1
X_15777_ game.CPU.applesa.ab.absxs.body_y\[105\] net446 vssd1 vssd1 vccd1 vccd1 _01789_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__12359__A game.CPU.applesa.ab.absxs.body_y\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19203__Q game.CPU.applesa.ab.XMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09647__B2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17516_ _02883_ _02915_ _02911_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11454__B2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12651__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14728_ _03505_ _08557_ vssd1 vssd1 vccd1 vccd1 _08560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_262_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18496_ net617 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__inv_2
XANTENNA__17185__A3 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19287__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12793__S net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17447_ net426 _02876_ _02833_ _02816_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__or4b_1
X_14659_ _04355_ _08490_ vssd1 vssd1 vccd1 vccd1 _08498_ sky130_fd_sc_hd__nor2_1
XFILLER_0_172_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09668__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17378_ net1119 net1121 _02806_ _02807_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14293__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19117_ net1182 _00157_ _00788_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[162\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16329_ net211 _02321_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__nand2_8
XFILLER_0_42_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09387__B net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10607__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16696__A2 _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19048_ net1186 _00280_ _00719_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[93\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_140_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_313_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13918__A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_301_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10717__B1 _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_336_Right_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16013__B net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13129__S net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13667__C1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ net912 game.CPU.applesa.ab.check_walls.above.walls\[56\] game.CPU.applesa.ab.check_walls.above.walls\[58\]
+ net922 _03945_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a221o_1
XFILLER_0_214_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11157__B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15852__B net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12968__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09886__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_A _06209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_241_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09634_ net1148 game.CPU.applesa.ab.absxs.body_y\[17\] vssd1 vssd1 vccd1 vccd1 _03877_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09850__B game.CPU.applesa.ab.absxs.body_y\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10996__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09565_ net1081 game.CPU.applesa.ab.absxs.body_x\[79\] vssd1 vssd1 vccd1 vccd1 _03808_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__09638__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09638__B2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11445__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12642__B1 game.CPU.applesa.twoapples.absxs.next_head\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09496_ net1130 net818 vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_322_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout807_A game.CPU.applesa.ab.check_walls.above.walls\[92\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_X net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_351_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_191_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18654__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_322_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09297__B game.CPU.applesa.ab.check_walls.above.walls\[81\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1337_X net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14147__B1 _07895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16687__A2 _02280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10340_ game.CPU.randy.f1.a1.count\[3\] net740 _04488_ game.CPU.randy.f1.a1.count\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_230_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19586__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10271_ game.CPU.applesa.ab.apple_possible\[4\] game.CPU.applesa.ab.apple_possible\[5\]
+ game.CPU.applesa.ab.apple_possible\[6\] game.CPU.applesa.ab.apple_possible\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__or4_1
XFILLER_0_103_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ _05332_ _05333_ _05336_ _05338_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__or4_1
XFILLER_0_264_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_303_Right_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15647__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12451__B net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_306_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout76_X net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout450 net451 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09463__D net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout461 net464 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__buf_2
Xfanout472 net475 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15762__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13961_ net867 net784 game.CPU.applesa.ab.check_walls.above.walls\[179\] net876 vssd1
+ vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11067__B net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout483 net486 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_2
Xfanout494 _06596_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_2
X_12912_ _06659_ _06660_ net692 vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__mux2_1
X_15700_ _01704_ _01705_ _01709_ _01710_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__or4b_1
X_16680_ net155 net100 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__nor2_1
XANTENNA__10487__A2 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11778__A1_N net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13892_ _07757_ _07758_ _07760_ _07765_ vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__or4_2
XFILLER_0_216_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12843_ game.writer.tracker.frame\[278\] game.writer.tracker.frame\[279\] net1018
+ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__mux2_1
X_15631_ net781 net431 net342 _03481_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__19023__Q game.CPU.applesa.ab.check_walls.above.walls\[68\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12859__S1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15562_ game.writer.updater.commands.mode\[2\] _06545_ _01580_ vssd1 vssd1 vccd1
+ vccd1 _01581_ sky130_fd_sc_hd__and3_1
XANTENNA__16086__A2_N net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18350_ net594 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__inv_2
XANTENNA__11436__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ _06644_ _06645_ _06647_ _06646_ net493 net686 vssd1 vssd1 vccd1 vccd1 _06648_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_83_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12633__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13830__C1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_291_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ net136 net114 _02379_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__or3b_1
XFILLER_0_28_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ game.CPU.apple_location2\[2\] net1053 vssd1 vssd1 vccd1 vccd1 _08387_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11725_ net573 _05338_ _05612_ _05333_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__o211a_1
X_15493_ _08926_ _01516_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__nand2_1
X_18281_ net622 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XFILLER_0_355_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13808__S0 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17232_ _02545_ net72 net730 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__o21a_1
XFILLER_0_327_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09488__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14444_ game.CPU.applesa.ab.absxs.body_y\[88\] net983 vssd1 vssd1 vccd1 vccd1 _08318_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__14386__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11656_ net829 net261 vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_155_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_330_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout90 net91 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_4
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17163_ net149 _02454_ net77 _02721_ net1513 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[452\]
+ sky130_fd_sc_hd__a32o_1
X_10607_ net1078 _04673_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__nor2_2
XANTENNA__11530__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14375_ game.CPU.applesa.ab.absxs.body_x\[118\] net879 net871 game.CPU.applesa.ab.absxs.body_y\[116\]
+ _08248_ vssd1 vssd1 vccd1 vccd1 _08249_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15002__B net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ game.CPU.applesa.ab.check_walls.above.walls\[107\] net762 vssd1 vssd1 vccd1
+ vccd1 _05476_ sky130_fd_sc_hd__xor2_2
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09801__B2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16114_ net446 game.CPU.applesa.ab.absxs.body_y\[69\] _03237_ net344 vssd1 vssd1
+ vccd1 vccd1 _02126_ sky130_fd_sc_hd__a2bb2o_1
X_13326_ _06730_ _06731_ _06740_ _06732_ net695 net480 vssd1 vssd1 vccd1 vccd1 _07200_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_134_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17094_ _02237_ net140 net560 vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10538_ game.CPU.applesa.ab.absxs.body_x\[44\] _04640_ _04641_ game.CPU.applesa.ab.absxs.body_x\[40\]
+ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__a22o_1
X_16045_ _03242_ net344 net334 _03309_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13257_ game.writer.tracker.frame\[452\] game.writer.tracker.frame\[453\] net1014
+ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__mux2_1
X_10469_ net1121 net1124 vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__nand2b_2
XANTENNA__09935__B net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12208_ game.CPU.applesa.ab.check_walls.above.walls\[142\] net417 vssd1 vssd1 vccd1
+ vccd1 _06094_ sky130_fd_sc_hd__xnor2_1
X_13188_ game.writer.tracker.frame\[438\] game.writer.tracker.frame\[439\] net1039
+ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_244_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12361__B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19804_ clknet_leaf_33_clk game.writer.tracker.next_frame\[399\] net1324 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[399\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11911__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15953__A game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _06021_ _06022_ _06023_ _06025_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__or4_2
X_17996_ net656 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__inv_2
XANTENNA__13113__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09951__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_341_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19735_ clknet_leaf_18_clk game.writer.tracker.next_frame\[330\] net1288 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[330\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15672__B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12788__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16947_ _02391_ net92 _02654_ net1491 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[302\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14569__A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11675__A1 game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19666_ clknet_leaf_29_clk game.writer.tracker.next_frame\[261\] net1291 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[261\] sky130_fd_sc_hd__dfrtp_1
X_16878_ _06703_ net148 _02298_ _02399_ net717 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__o41a_1
XANTENNA__16602__A2 _02455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18617_ clknet_leaf_13_clk _01034_ _00354_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[111\]
+ sky130_fd_sc_hd__dfrtp_4
X_15829_ game.CPU.applesa.ab.absxs.body_x\[16\] net273 vssd1 vssd1 vccd1 vccd1 _01841_
+ sky130_fd_sc_hd__nand2_1
X_19597_ clknet_leaf_35_clk game.writer.tracker.next_frame\[192\] net1355 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[192\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_273_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12089__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_338_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09350_ _03588_ _03589_ _03590_ _03592_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__a211o_1
X_18548_ net626 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__inv_2
XANTENNA__18677__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19922__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_255_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18772__Q game.CPU.applesa.ab.absxs.body_x\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_318_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09281_ game.CPU.applesa.ab.check_walls.above.walls\[196\] game.CPU.applesa.ab.check_walls.above.walls\[197\]
+ game.CPU.applesa.ab.check_walls.above.walls\[198\] net780 vssd1 vssd1 vccd1 vccd1
+ _03526_ sky130_fd_sc_hd__nor4_1
XFILLER_0_129_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18479_ net635 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_177_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09398__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16008__B net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12536__B net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11440__B net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout123_A _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11562__A2_N net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_344_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload60 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__inv_16
Xclkload71 clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__inv_6
XFILLER_0_286_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_266_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout492_A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15629__B1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11902__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__A game.CPU.applesa.ab.absxs.body_y\[76\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15863__A game.CPU.applesa.ab.absxs.body_x\[114\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08996_ game.CPU.applesa.ab.absxs.body_x\[37\] vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__inv_2
XANTENNA__16678__B _02237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16841__A2 _02299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout280_X net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19452__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16054__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ net1140 game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1
+ vccd1 _03860_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_355_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout924_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_203_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11418__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09548_ net1132 game.CPU.applesa.ab.absxs.body_y\[115\] vssd1 vssd1 vccd1 vccd1 _03791_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_277_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12615__B1 _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18682__Q game.CPU.applesa.ab.absxs.body_x\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16357__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09479_ _03719_ _03720_ _03721_ _03718_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__a211o_1
XFILLER_0_182_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ game.CPU.applesa.ab.check_walls.above.walls\[3\] net764 vssd1 vssd1 vccd1
+ vccd1 _05399_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12490_ _03266_ game.CPU.applesa.twoapples.absxs.next_head\[0\] vssd1 vssd1 vccd1
+ vccd1 _06367_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10641__A2 game.CPU.applesa.ab.absxs.body_x\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12446__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12918__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11441_ net825 net261 _05329_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14160_ net926 net1048 net866 net1150 vssd1 vssd1 vccd1 vccd1 _08034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_278_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15757__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11372_ net568 _05254_ _05258_ _05259_ _05260_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__a2111o_1
XANTENNA__08940__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12733__Y _06607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13111_ game.writer.tracker.frame\[144\] game.writer.tracker.frame\[145\] net1023
+ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__mux2_2
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10323_ _04501_ _04502_ vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_308_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09755__B net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14091_ net1075 game.CPU.applesa.ab.check_walls.above.walls\[8\] vssd1 vssd1 vccd1
+ vccd1 _07965_ sky130_fd_sc_hd__xor2_1
XFILLER_0_277_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13042_ _06870_ _06885_ net697 vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__mux2_1
X_10254_ net759 net571 _04446_ net1173 vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_5_Left_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12181__B _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__buf_2
X_17850_ _01445_ _03174_ net182 vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__a21o_1
Xfanout1212 net1216 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__buf_2
X_10185_ _04363_ _04371_ _04374_ _04365_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__a31o_1
Xfanout1223 net1224 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16588__B net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1234 net1235 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__buf_1
X_16801_ _02485_ net104 _02601_ net1661 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[210\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_206_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1245 net1246 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__buf_1
XANTENNA__16832__A2 _02369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1256 net1257 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__clkbuf_2
X_17781_ net1991 _03125_ _03130_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__a21oi_1
Xfanout1267 game.CPU.applesa.ab.absxs.body_x\[76\] vssd1 vssd1 vccd1 vccd1 net1267
+ sky130_fd_sc_hd__buf_4
XANTENNA__13646__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout280 _06610_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_4
Xfanout1278 net26 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__buf_2
X_14993_ net1223 net1250 game.CPU.applesa.ab.check_walls.above.walls\[21\] vssd1 vssd1
+ vccd1 vccd1 _00209_ sky130_fd_sc_hd__and3_1
Xfanout291 net292 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_4
X_19520_ clknet_leaf_21_clk game.writer.tracker.next_frame\[115\] net1317 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[115\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13293__A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1289 net1290 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11806__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12854__A0 _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16732_ _02514_ net62 _02580_ net1544 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[162\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13944_ net870 game.CPU.applesa.ab.check_walls.above.walls\[68\] game.CPU.applesa.ab.check_walls.above.walls\[70\]
+ net854 _07813_ vssd1 vssd1 vccd1 vccd1 _07818_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16045__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19945__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19451_ clknet_leaf_49_clk game.writer.tracker.next_frame\[46\] net1295 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[46\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11525__B net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16663_ net168 net154 _02348_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__and3_1
XANTENNA__16596__A1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13875_ net960 game.CPU.applesa.ab.check_walls.above.walls\[109\] vssd1 vssd1 vccd1
+ vccd1 _07749_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_319_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18402_ net618 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__inv_2
X_12826_ _06633_ _06635_ _06637_ _06632_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__o31a_1
X_15614_ game.CPU.applesa.ab.check_walls.above.walls\[83\] net458 vssd1 vssd1 vccd1
+ vccd1 _01626_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12606__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19382_ clknet_leaf_3_clk _01388_ _00962_ vssd1 vssd1 vccd1 vccd1 game.CPU.bodymain1.main.score\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_16594_ _02351_ _02439_ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__nand2_1
XFILLER_0_347_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18333_ net594 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__inv_2
X_12757_ _06627_ _06628_ _06630_ _06629_ net476 net677 vssd1 vssd1 vccd1 vccd1 _06631_
+ sky130_fd_sc_hd__mux4_1
X_15545_ net954 _01545_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_315_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11708_ _05583_ _05595_ _05596_ _05582_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__o31a_1
XANTENNA__15013__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16899__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15476_ _08879_ _01467_ _01492_ _01501_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__a22o_1
XFILLER_0_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11290__C1 _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18264_ net649 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__inv_2
XFILLER_0_355_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12688_ net888 net879 vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__nor2_1
XFILLER_0_315_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12356__B net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12909__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17215_ _02299_ net142 net119 _02734_ net1789 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[491\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14427_ game.CPU.applesa.ab.absxs.body_x\[25\] net1061 vssd1 vssd1 vccd1 vccd1 _08301_
+ sky130_fd_sc_hd__xnor2_1
X_11639_ game.CPU.applesa.ab.check_walls.above.walls\[152\] net774 vssd1 vssd1 vccd1
+ vccd1 _05528_ sky130_fd_sc_hd__xnor2_1
X_18195_ net608 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__inv_2
XFILLER_0_330_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18324__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13582__A1 game.writer.tracker.frame\[375\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19325__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17146_ _02419_ net58 net560 vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_250_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14358_ game.CPU.applesa.ab.absxs.body_y\[103\] net941 vssd1 vssd1 vccd1 vccd1 _08232_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_3_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_268_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13309_ net504 _06758_ net699 vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17077_ _02464_ net60 _02695_ net2022 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[392\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_268_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16520__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_268_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12372__A game.CPU.applesa.ab.absxs.body_x\[114\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14289_ _08160_ _08161_ _08162_ vssd1 vssd1 vccd1 vccd1 _08163_ sky130_fd_sc_hd__and3_1
XANTENNA__09665__B game.CPU.applesa.ab.absxs.body_y\[38\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13334__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14531__B1 _07742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16028_ _03297_ net340 net432 game.CPU.applesa.ab.absxs.body_y\[95\] vssd1 vssd1
+ vccd1 vccd1 _02040_ sky130_fd_sc_hd__a22o_1
XANTENNA__12091__B net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19475__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17076__A2 _02373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10699__A2 _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13915__B game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17979_ net605 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__inv_2
XFILLER_0_354_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13407__S net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19718_ clknet_leaf_35_clk game.writer.tracker.next_frame\[313\] net1345 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[313\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09710__B1 game.CPU.applesa.ab.absxs.body_y\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19649_ clknet_leaf_21_clk game.writer.tracker.next_frame\[244\] net1337 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[244\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16587__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09402_ net895 net807 net805 net904 _03643_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__a221o_1
XFILLER_0_177_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13931__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09333_ _03572_ _03573_ _03574_ _03575_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout240_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17000__A2 _02670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_303_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10623__A2 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09264_ game.CPU.randy.counter1.count\[3\] vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11820__A1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_350_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11820__B2 game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12266__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11170__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09195_ game.CPU.applesa.ab.check_walls.above.walls\[121\] vssd1 vssd1 vccd1 vccd1
+ _03444_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout126_X net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout505_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1247_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09856__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_214_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15577__B net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11584__B1 _05408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19818__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12282__A game.CPU.applesa.ab.check_walls.above.walls\[133\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13325__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09529__B1 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17792__B net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_328_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1202_X net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 game.CPU.right_button.eD1.D vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_328_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold22 game.CPU.left_button.eD1.Q1 vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16814__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold33 game.CPU.applesa.normal1.number\[3\] vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_303_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold44 game.CPU.applesa.twomode.number\[6\] vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ game.CPU.applesa.ab.absxs.body_x\[95\] vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__inv_2
XFILLER_0_264_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold55 net48 vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_279_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11626__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold66 game.CPU.applesa.ab.absxs.body_y\[0\] vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12836__A0 game.writer.tracker.frame\[320\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold77 game.CPU.applesa.steady\[0\] vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 game.writer.tracker.frame\[246\] vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14002__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11990_ _05320_ _05321_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__nand2_1
Xhold99 game.writer.tracker.frame\[442\] vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ _04827_ _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout927_X net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09482__A1_N net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13660_ _07532_ _07533_ net481 vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__mux2_1
X_10872_ game.CPU.randy.counter1.count\[18\] _03495_ _04766_ _04774_ vssd1 vssd1 vccd1
+ vccd1 game.CPU.randy.counter1.out sky130_fd_sc_hd__o22a_2
XTAP_TAPCELL_ROW_67_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_356_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19948__RESET_B net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12611_ game.CPU.applesa.ab.absxs.body_y\[21\] net526 net363 game.CPU.applesa.ab.absxs.body_y\[20\]
+ _06424_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__o221a_1
XFILLER_0_168_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12064__A1 game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13591_ game.writer.tracker.frame\[349\] game.writer.tracker.frame\[351\] game.writer.tracker.frame\[352\]
+ game.writer.tracker.frame\[350\] net975 net1017 vssd1 vssd1 vccd1 vccd1 _07465_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12064__B2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_197_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15330_ game.CPU.applesa.twomode.number\[7\] _08870_ vssd1 vssd1 vccd1 vccd1 _08873_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11361__A game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19348__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12542_ game.CPU.applesa.ab.absxs.body_x\[41\] net380 game.CPU.applesa.twoapples.absxs.next_head\[4\]
+ _03344_ _06418_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__a221o_1
XANTENNA__10614__A2 _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_314_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13239__S1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15261_ game.CPU.kyle.L1.nextState\[1\] _08809_ _08810_ net1871 vssd1 vssd1 vccd1
+ vccd1 _08818_ sky130_fd_sc_hd__a22oi_4
X_12473_ game.CPU.applesa.ab.absxs.body_x\[56\] net382 vssd1 vssd1 vccd1 vccd1 _06350_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_152_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16750__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17000_ _02322_ _02670_ net729 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14212_ game.CPU.applesa.ab.absxs.body_y\[92\] net983 vssd1 vssd1 vccd1 vccd1 _08086_
+ sky130_fd_sc_hd__or2_1
XANTENNA__13564__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ _05296_ _05299_ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__and3_1
XFILLER_0_340_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15192_ _08760_ _08763_ game.CPU.walls.enable_in2 _08754_ vssd1 vssd1 vccd1 vccd1
+ _00016_ sky130_fd_sc_hd__o211ai_2
XANTENNA__19498__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_8 _02179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _08000_ _08003_ _08016_ _07916_ _07745_ vssd1 vssd1 vccd1 vccd1 _08017_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_340_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11355_ game.CPU.applesa.ab.check_walls.above.walls\[141\] net314 vssd1 vssd1 vccd1
+ vccd1 _05244_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_78_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13316__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_238_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ game.CPU.randy.f1.a1.count\[4\] game.CPU.randy.f1.a1.count\[3\] _04488_ vssd1
+ vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__and3_1
X_14074_ net870 net832 game.CPU.applesa.ab.check_walls.above.walls\[6\] net853 vssd1
+ vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__o22a_1
X_18951_ clknet_leaf_67_clk net1406 _00622_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11286_ _04984_ _04986_ _04987_ _04988_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16599__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13867__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17058__A2 _02670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13025_ _06897_ _06898_ net485 vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__mux2_1
X_17902_ net661 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__inv_2
XFILLER_0_238_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11878__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10237_ _04395_ _04398_ _04397_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__a21oi_1
X_18882_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[12\] _00577_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[12\] sky130_fd_sc_hd__dfrtp_1
Xfanout1020 net1022 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_4
Xfanout1031 net1034 vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_238_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16805__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17833_ _03161_ _03162_ game.writer.updater.commands.count\[5\] net182 vssd1 vssd1
+ vccd1 vccd1 _01414_ sky130_fd_sc_hd__a2bb2o_1
Xfanout1042 game.CPU.applesa.y\[0\] vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_218_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1053 net1054 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__clkbuf_8
X_10168_ game.CPU.randy.f1.c1.max_i\[0\] _04341_ _04361_ vssd1 vssd1 vccd1 vccd1 _01334_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_163_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10550__A1 game.CPU.applesa.ab.absxs.body_x\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10550__B2 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1064 net1068 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13227__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1075 net1077 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__buf_6
XANTENNA__11536__A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1086 net1087 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__buf_4
XANTENNA__15008__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17764_ game.CPU.applesa.twoapples.count_luck\[4\] _03116_ vssd1 vssd1 vccd1 vccd1
+ _03119_ sky130_fd_sc_hd__nand2_1
Xfanout1097 net1099 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__buf_4
XFILLER_0_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14976_ net1225 net1252 net832 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__and3_1
X_10099_ _04298_ _04301_ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__or3b_1
XFILLER_0_107_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19503_ clknet_leaf_26_clk game.writer.tracker.next_frame\[98\] net1313 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[98\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_261_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16715_ net185 _02498_ net106 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__and3_1
XFILLER_0_348_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13927_ net1055 game.CPU.applesa.ab.check_walls.above.walls\[34\] vssd1 vssd1 vccd1
+ vccd1 _07801_ sky130_fd_sc_hd__xor2_1
X_17695_ game.CPU.walls.rand_wall.input2 net580 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_347_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19434_ clknet_leaf_39_clk game.writer.tracker.next_frame\[29\] net1352 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[29\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17230__A2 _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16646_ _02407_ _02520_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_179_Right_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13858_ game.writer.tracker.frame\[557\] game.writer.tracker.frame\[559\] game.writer.tracker.frame\[560\]
+ game.writer.tracker.frame\[558\] net972 net1007 vssd1 vssd1 vccd1 vccd1 _07732_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_186_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14566__B _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_347_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12809_ game.writer.tracker.frame\[364\] game.writer.tracker.frame\[365\] net998
+ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19365_ clknet_leaf_69_clk _01371_ _00946_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16577_ net150 net126 _02498_ _02495_ net1747 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[89\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_44_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19211__Q game.CPU.applesa.ab.apple_possible\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13789_ _07661_ _07662_ net496 vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_252_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19618__RESET_B net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18316_ net615 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15528_ net1049 _01549_ _06557_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__mux2_1
XANTENNA__10605__A2 _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_328_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19296_ clknet_leaf_69_clk net326 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.x_final\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18715__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18247_ net645 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
XANTENNA__16741__A1 _02378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15459_ _01456_ _01481_ _01483_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_316_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09676__A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18178_ net608 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13198__A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold503 game.writer.tracker.frame\[53\] vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_68_Left_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_279_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17129_ net165 _02386_ net76 _02711_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[428\]
+ sky130_fd_sc_hd__a31o_1
Xhold514 game.writer.updater.commands.count\[1\] vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17893__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold525 game.CPU.randy.f1.a1.count\[10\] vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 game.writer.tracker.frame\[533\] vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 game.writer.tracker.frame\[2\] vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 game.writer.tracker.frame\[556\] vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14504__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ net1119 _04175_ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_284_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold569 game.writer.tracker.frame\[528\] vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload25_A clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_263_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17049__A2 _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13926__A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09882_ _03792_ _03794_ _03796_ _03930_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__o31a_2
XANTENNA__11869__A1 _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16302__A _06573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12530__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout190_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_224_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16021__B net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13137__S net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout288_A net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10541__B2 game.CPU.applesa.ab.absxs.body_x\[35\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14283__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Left_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15860__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_352_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1197_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17221__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_314_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_274_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16980__A1 _02458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout243_X net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout622_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11181__A game.CPU.applesa.ab.absxs.body_x\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_353_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_216_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09316_ net1140 game.CPU.applesa.ab.absxs.body_y\[66\] vssd1 vssd1 vccd1 vccd1 _03559_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__13794__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18960__Q game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09247_ game.CPU.randy.counter1.count1\[18\] vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__inv_2
XFILLER_0_330_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19640__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16732__A1 _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1152_X net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13600__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12349__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13546__B2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09586__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09178_ game.CPU.applesa.ab.check_walls.above.walls\[88\] vssd1 vssd1 vccd1 vccd1
+ _03427_ sky130_fd_sc_hd__inv_2
XFILLER_0_279_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout991_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12724__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14412__A1_N game.CPU.applesa.ab.absxs.body_x\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17288__A2 _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_322_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput12 net12 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
X_11140_ _05022_ _05023_ _05025_ _05026_ _05028_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_9_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XANTENNA__19790__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_285_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13849__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_101_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_227_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11071_ _04952_ _04953_ _04956_ _04957_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a211o_1
XFILLER_0_290_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_275_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10022_ _04225_ _04228_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__nand2b_1
XANTENNA__16799__A1 _02483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19020__CLK net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16799__B2 game.writer.tracker.frame\[209\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__A game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14830_ game.CPU.randy.f1.c1.count\[0\] game.CPU.randy.f1.c1.count\[1\] game.CPU.randy.f1.c1.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _08632_ sky130_fd_sc_hd__and3_1
XFILLER_0_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14274__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15770__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11075__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__S net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14761_ game.CPU.randy.counter1.count\[15\] net265 _08581_ game.CPU.randy.counter1.count\[13\]
+ vssd1 vssd1 vccd1 vccd1 _08582_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11973_ game.CPU.applesa.ab.apple_possible\[6\] _05192_ vssd1 vssd1 vccd1 vccd1 _05860_
+ sky130_fd_sc_hd__nand2_1
X_16500_ net154 _02444_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_329_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13712_ game.writer.tracker.frame\[205\] game.writer.tracker.frame\[207\] game.writer.tracker.frame\[208\]
+ game.writer.tracker.frame\[206\] net974 net1010 vssd1 vssd1 vccd1 vccd1 _07586_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__17212__A2 _02720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10924_ net541 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.next_head\[6\] sky130_fd_sc_hd__inv_2
XANTENNA__19170__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17480_ _02902_ _02908_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__nand2_1
X_14692_ game.CPU.randy.counter1.count1\[13\] _08500_ _08530_ game.CPU.randy.counter1.count1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _08531_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_316_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13234__A0 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16431_ _02350_ _02372_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__or2_2
XFILLER_0_128_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_345_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13643_ game.writer.tracker.frame\[31\] net711 net674 game.writer.tracker.frame\[32\]
+ vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__o22a_1
XANTENNA__18738__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12037__B2 game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17978__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11803__B net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855_ _03498_ game.CPU.randy.counter1.count1\[15\] _03499_ game.CPU.randy.counter1.count1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a22o_1
XANTENNA__16971__A1 _02436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_238_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12187__A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16882__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16971__B2 game.writer.tracker.frame\[320\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_317_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13785__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_clk_X clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19150_ net1188 _00193_ _00821_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[195\]
+ sky130_fd_sc_hd__dfrtp_4
X_16362_ _02343_ _02345_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__or2_1
X_13574_ _07446_ _07447_ net502 vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__mux2_1
X_10786_ net932 game.CPU.applesa.ab.absxs.body_y\[47\] net562 _04724_ vssd1 vssd1
+ vccd1 vccd1 _01006_ sky130_fd_sc_hd__a31o_1
XFILLER_0_109_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18101_ net603 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__inv_2
XANTENNA__10419__B _04563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15313_ game.CPU.applesa.twomode.number\[4\] _08854_ vssd1 vssd1 vccd1 vccd1 _08859_
+ sky130_fd_sc_hd__or2_1
X_12525_ game.CPU.applesa.ab.absxs.body_x\[96\] net381 vssd1 vssd1 vccd1 vccd1 _06402_
+ sky130_fd_sc_hd__or2_1
X_16293_ game.writer.tracker.frame\[11\] net720 _02292_ vssd1 vssd1 vccd1 vccd1 _02293_
+ sky130_fd_sc_hd__and3_1
X_19081_ net1186 _00117_ _00752_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16723__A1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_240_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15526__A2 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16184__C1 _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18032_ net589 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__inv_2
XANTENNA__18888__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09496__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15244_ game.CPU.kyle.L1.cnt_500hz\[13\] game.CPU.kyle.L1.cnt_500hz\[14\] game.CPU.kyle.L1.cnt_500hz\[12\]
+ vssd1 vssd1 vccd1 vccd1 _08805_ sky130_fd_sc_hd__and3b_1
X_12456_ net1269 net380 net526 game.CPU.applesa.ab.absxs.body_y\[49\] vssd1 vssd1
+ vccd1 vccd1 _06333_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_240_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11548__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11407_ net797 net255 vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__nand2_1
XANTENNA__17279__A2 _02574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15175_ _04582_ _04584_ _08749_ net1116 vssd1 vssd1 vccd1 vccd1 _08751_ sky130_fd_sc_hd__a211o_1
XANTENNA__15010__B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12387_ game.CPU.applesa.ab.absxs.body_y\[24\] net363 vssd1 vssd1 vccd1 vccd1 _06264_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_327_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_297_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14126_ net1065 _03391_ game.CPU.applesa.ab.check_walls.above.walls\[28\] net870
+ _07995_ vssd1 vssd1 vccd1 vccd1 _08000_ sky130_fd_sc_hd__o221a_1
XFILLER_0_249_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11338_ game.CPU.applesa.ab.check_walls.above.walls\[81\] net770 vssd1 vssd1 vccd1
+ vccd1 _05227_ sky130_fd_sc_hd__xor2_1
XFILLER_0_278_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19983_ clknet_leaf_46_clk _01407_ net1280 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.y\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_265_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10771__B2 game.CPU.applesa.ab.absxs.body_y\[69\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13746__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18934_ clknet_leaf_14_clk net1398 net1282 vssd1 vssd1 vccd1 vccd1 game.CPU.reset_button1.eD1.Q1
+ sky130_fd_sc_hd__dfrtp_1
X_14057_ net948 game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1 vccd1
+ vccd1 _07931_ sky130_fd_sc_hd__xor2_1
X_11269_ _05014_ _05015_ _05017_ _05018_ _05147_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_248_Right_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15647__A2_N net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13008_ game.writer.tracker.frame\[560\] game.writer.tracker.frame\[561\] net1007
+ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__mux2_1
XANTENNA__12512__A2 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18865_ clknet_leaf_0_clk _01256_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_253_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14273__A2_N net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19206__Q game.CPU.applesa.ab.YMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17816_ _08894_ net576 _01438_ _01444_ _03147_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__o221a_2
XFILLER_0_175_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10170__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17451__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18796_ clknet_leaf_4_clk _00039_ _00533_ vssd1 vssd1 vccd1 vccd1 game.CPU.bodymain1.main.pause_clk
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__19513__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14265__A2 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_261_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15680__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17747_ net757 game.CPU.applesa.twomode.counter_normal vssd1 vssd1 vccd1 vccd1 _01348_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__11079__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14959_ _08672_ _08674_ _08667_ _08671_ vssd1 vssd1 vccd1 vccd1 _08736_ sky130_fd_sc_hd__o211a_1
XANTENNA__18049__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_342_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_338_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17203__A2 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17678_ game.CPU.walls.rand_wall.count_luck\[1\] _03063_ vssd1 vssd1 vccd1 vccd1
+ _03065_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16411__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14296__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13225__A0 _07096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19417_ clknet_leaf_48_clk game.writer.tracker.next_frame\[12\] net1303 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16629_ net1764 _02532_ _02533_ net124 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[106\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11713__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17888__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16962__A1 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19663__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13776__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19348_ clknet_leaf_70_clk game.CPU.applesa.twoapples.absxs.next_head\[4\] vssd1
+ vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.y_final\[0\] sky130_fd_sc_hd__dfxtp_1
X_09101_ game.CPU.applesa.ab.absxs.body_y\[25\] vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__inv_2
XFILLER_0_162_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16714__A1 _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19279_ clknet_leaf_65_clk game.CPU.applesa.ab.absxs.collision vssd1 vssd1 vccd1
+ vccd1 game.CPU.applesa.ab.collisions sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13420__S net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09032_ game.CPU.applesa.ab.absxs.body_x\[24\] vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12544__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16016__B net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold300 game.writer.tracker.frame\[347\] vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_304_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_211_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold311 game.writer.tracker.frame\[400\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_276_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout203_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 game.writer.tracker.frame\[77\] vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18512__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16478__B1 _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold333 game.writer.tracker.frame\[498\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 game.writer.tracker.frame\[367\] vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 game.writer.tracker.frame\[183\] vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold366 _04322_ vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 game.writer.tracker.frame\[194\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 game.writer.tracker.frame\[335\] vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_6_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout802 game.CPU.applesa.ab.check_walls.above.walls\[103\] vssd1 vssd1 vccd1 vccd1
+ net802 sky130_fd_sc_hd__clkbuf_4
Xhold399 game.writer.tracker.frame\[322\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_272_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09934_ game.CPU.bodymain1.main.score\[0\] _03527_ _04158_ vssd1 vssd1 vccd1 vccd1
+ _04172_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1112_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout813 game.CPU.applesa.ab.check_walls.above.walls\[77\] vssd1 vssd1 vccd1 vccd1
+ net813 sky130_fd_sc_hd__clkbuf_4
Xfanout824 game.CPU.applesa.ab.check_walls.above.walls\[36\] vssd1 vssd1 vccd1 vccd1
+ net824 sky130_fd_sc_hd__clkbuf_4
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_215_Right_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10999__B net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_271_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout846 _04253_ vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__buf_4
XANTENNA__09904__B1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20054_ net1372 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
X_09865_ _04098_ _04099_ _04105_ _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__a211o_1
Xfanout857 _03376_ vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__buf_4
XANTENNA_input8_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10514__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout572_A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout868 _03374_ vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_4
Xfanout879 net880 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09380__A1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09380__B2 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_300_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ net916 game.CPU.applesa.ab.absxs.body_x\[41\] _03344_ net1158 vssd1 vssd1
+ vccd1 vccd1 _04039_ sky130_fd_sc_hd__o22a_1
XANTENNA__18955__Q game.CPU.applesa.ab.check_walls.above.walls\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_222_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14487__A _08053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10817__A2 game.CPU.applesa.ab.absxs.body_y\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09683__A2 game.CPU.applesa.ab.absxs.body_y\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12719__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_327_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11623__B net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16953__A1 _02404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10640_ _03273_ net561 vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_194_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10571_ _04580_ _04591_ _04617_ _04595_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a31o_2
XANTENNA__12294__X _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16705__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12735__A _06607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_311_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12310_ game.CPU.applesa.ab.check_walls.above.walls\[191\] net421 vssd1 vssd1 vccd1
+ vccd1 _06196_ sky130_fd_sc_hd__or2_1
XFILLER_0_334_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13290_ _06859_ _06922_ _07163_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__or3_2
XFILLER_0_16_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout994_X net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__Y _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12241_ game.CPU.applesa.ab.check_walls.above.walls\[151\] net422 vssd1 vssd1 vccd1
+ vccd1 _06127_ sky130_fd_sc_hd__nor2_1
XFILLER_0_267_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16469__B1 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12172_ _05282_ _05283_ _05284_ _05286_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__or4b_2
XANTENNA__15765__B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10753__B2 game.CPU.applesa.ab.absxs.body_y\[106\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11123_ game.CPU.applesa.ab.absxs.body_y\[18\] net401 vssd1 vssd1 vccd1 vccd1 _05013_
+ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09763__B game.CPU.applesa.ab.check_walls.above.walls\[98\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16980_ _02458_ net90 _02665_ net1944 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[325\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19536__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11054_ game.CPU.applesa.ab.absxs.body_y\[107\] net398 vssd1 vssd1 vccd1 vccd1 _04944_
+ sky130_fd_sc_hd__xnor2_1
X_15931_ game.CPU.applesa.ab.check_walls.above.walls\[127\] net430 vssd1 vssd1 vccd1
+ vccd1 _01943_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19026__Q game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10505__A1 net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_322_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10505__B2 game.CPU.applesa.ab.absxs.body_x\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10005_ net1105 _04212_ _04211_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09371__A1 net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18650_ clknet_leaf_51_clk _01067_ _00387_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[60\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09371__B2 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15862_ game.CPU.applesa.ab.absxs.body_x\[112\] net355 vssd1 vssd1 vccd1 vccd1 _01874_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__19963__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17601_ _03003_ _03016_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_58_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14813_ _08621_ _08622_ vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__nor2_1
X_18581_ clknet_leaf_53_clk _01001_ _00318_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[42\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__18560__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15793_ net1269 net352 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19686__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15995__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13550__S0 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17532_ _02948_ _02953_ _02959_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__or3_1
XANTENNA__11814__A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14744_ net55 _08569_ _08570_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__and3_1
XANTENNA__10808__A2 _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11956_ game.CPU.applesa.ab.check_walls.above.walls\[71\] net311 vssd1 vssd1 vccd1
+ vccd1 _05844_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_86_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14304__A1_N game.CPU.applesa.ab.absxs.body_y\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_357_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10907_ net1273 game.CPU.luck1.Qa\[0\] _04733_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__mux2_1
X_17463_ _02887_ _02888_ _02889_ _02791_ _08750_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__o32a_1
XANTENNA__15005__B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11887_ game.CPU.applesa.ab.check_walls.above.walls\[20\] net393 vssd1 vssd1 vccd1
+ vccd1 _05775_ sky130_fd_sc_hd__nand2_1
X_14675_ game.CPU.randy.counter1.count1\[3\] _04356_ vssd1 vssd1 vccd1 vccd1 _08514_
+ sky130_fd_sc_hd__and2_1
X_19202_ clknet_leaf_67_clk net1435 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16414_ net115 net159 _02382_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13626_ game.writer.tracker.frame\[309\] game.writer.tracker.frame\[311\] game.writer.tracker.frame\[312\]
+ game.writer.tracker.frame\[310\] net979 net1033 vssd1 vssd1 vccd1 vccd1 _07500_
+ sky130_fd_sc_hd__mux4_1
X_10838_ game.CPU.randy.counter1.count\[11\] _03502_ _03503_ game.CPU.randy.counter1.count1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_27_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17394_ _04808_ _02778_ _02818_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__and3b_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_305_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_333_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12966__C1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19133_ net1183 _00174_ _00804_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[178\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_333_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16345_ net1971 net732 _02329_ _02332_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[23\]
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12430__A1 net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13557_ game.writer.tracker.frame\[102\] net841 net709 game.writer.tracker.frame\[103\]
+ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__o22a_1
XFILLER_0_109_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10769_ game.CPU.applesa.ab.absxs.body_y\[75\] _04675_ _04676_ game.CPU.applesa.ab.absxs.body_y\[71\]
+ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12430__B2 game.CPU.applesa.ab.absxs.body_x\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_332_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_317_Right_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19064_ net1186 _00098_ _00735_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[109\]
+ sky130_fd_sc_hd__dfrtp_4
X_12508_ game.CPU.applesa.ab.absxs.body_y\[75\] net367 vssd1 vssd1 vccd1 vccd1 _06385_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_298_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13488_ net209 _07358_ _07361_ net284 vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__a211o_1
X_16276_ net134 net70 _02280_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_11_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_298_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16172__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19066__CLK net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18015_ net657 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__inv_2
XFILLER_0_258_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15956__A game.CPU.applesa.ab.check_walls.above.walls\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12439_ game.CPU.applesa.ab.absxs.body_x\[104\] net382 vssd1 vssd1 vccd1 vccd1 _06316_
+ sky130_fd_sc_hd__or2_1
X_15227_ game.CPU.applesa.normal1.counter _08788_ _08789_ _08790_ _08791_ vssd1 vssd1
+ vccd1 vccd1 _08792_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10165__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16404__X _02375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12733__A2 _06571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17121__A1 _02370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15675__B net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15158_ net1213 net1240 game.CPU.applesa.ab.check_walls.above.walls\[186\] vssd1
+ vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__and3_1
XFILLER_0_238_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_247_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_292_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14109_ _07975_ _07981_ _07982_ vssd1 vssd1 vccd1 vccd1 _07983_ sky130_fd_sc_hd__and3_1
Xfanout109 net110 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__clkbuf_4
X_19966_ clknet_leaf_41_clk game.writer.tracker.next_frame\[561\] net1327 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[561\] sky130_fd_sc_hd__dfrtp_1
X_15089_ net1206 net1232 net798 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__and3_1
XFILLER_0_266_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18917_ clknet_leaf_5_clk net1394 _00601_ vssd1 vssd1 vccd1 vccd1 game.CPU.up_button.eD1.D
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19897_ clknet_leaf_15_clk game.writer.tracker.next_frame\[492\] net1293 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[492\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_219_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09898__C1 _04140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18903__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09650_ net1145 game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1 vssd1 vccd1
+ vccd1 _03893_ sky130_fd_sc_hd__xor2_1
XANTENNA__15691__A game.CPU.applesa.ab.absxs.body_y\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_241_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18848_ clknet_leaf_0_clk _01239_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_124_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09581_ net916 game.CPU.applesa.ab.check_walls.above.walls\[41\] game.CPU.applesa.ab.check_walls.above.walls\[45\]
+ net900 _03817_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__a221o_1
X_18779_ clknet_leaf_63_clk _01196_ _00516_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[93\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_261_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13541__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17188__A1 _02494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14100__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17114__C net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_258_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11443__B net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11472__A2 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout153_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16935__A1 _02370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18507__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_271_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17411__A net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10680__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12957__C1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19409__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12421__A1 game.CPU.applesa.ab.absxs.body_x\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout320_A game.CPU.applesa.ab.absxs.next_head\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12421__B2 game.CPU.applesa.ab.absxs.body_x\[35\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout418_A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1062_A game.CPU.applesa.x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_311_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_304_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12274__B net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09015_ game.CPU.applesa.ab.absxs.body_x\[88\] vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14174__B2 game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout206_X net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18242__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19559__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1327_A net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 game.writer.tracker.frame\[321\] vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13921__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 game.writer.tracker.frame\[206\] vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13921__B2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17112__A1 _02359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_269_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold152 game.writer.tracker.frame\[292\] vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 game.writer.tracker.frame\[314\] vssd1 vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__B2 game.CPU.applesa.ab.absxs.body_y\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold174 game.writer.tracker.frame\[454\] vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 game.writer.tracker.frame\[178\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09583__B net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_282_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold196 game.writer.tracker.frame\[403\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 net612 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_4
XANTENNA__14477__A2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout621 net623 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_224_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11618__B net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09917_ net930 _04156_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__nand2_2
Xfanout632 net633 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_298_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout643 net646 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__buf_4
XANTENNA_fanout954_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout654 net655 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_4
XANTENNA__18583__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_X net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout665 net667 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__buf_4
XANTENNA__09353__A1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout676 net677 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__buf_4
XFILLER_0_336_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20037_ net1385 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XANTENNA__09353__B2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout687 net691 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_4
X_09848_ net925 game.CPU.applesa.ab.absxs.body_x\[31\] game.CPU.applesa.ab.absxs.body_y\[31\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__a22o_1
Xfanout698 net699 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_109_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_336_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18685__Q game.CPU.applesa.ab.absxs.body_x\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_225_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_358_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09779_ net1127 net789 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_358_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ game.CPU.applesa.ab.check_walls.above.walls\[62\] net302 _05691_ _05692_
+ _05697_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__o2111a_1
XANTENNA__13988__A1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12790_ game.writer.tracker.frame\[382\] game.writer.tracker.frame\[383\] net1032
+ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_240_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13988__B2 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12449__B game.CPU.applesa.twoapples.absxs.next_head\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11999__B1 _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__B net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ _04441_ _05524_ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09104__A game.CPU.applesa.ab.absxs.body_y\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16926__A1 _02434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_235_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _08331_ _08332_ _08333_ _08326_ vssd1 vssd1 vccd1 vccd1 _08334_ sky130_fd_sc_hd__a211o_1
X_11672_ game.CPU.applesa.ab.check_walls.above.walls\[127\] net258 vssd1 vssd1 vccd1
+ vccd1 _05561_ sky130_fd_sc_hd__nand2_1
XANTENNA__08943__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14401__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12948__C1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_315_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13411_ net680 _06875_ _07284_ net507 vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__o211a_1
X_10623_ game.CPU.applesa.ab.absxs.body_x\[66\] _04679_ _04680_ game.CPU.applesa.ab.absxs.body_x\[62\]
+ vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12412__A1 game.CPU.applesa.ab.absxs.body_x\[55\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14391_ game.CPU.applesa.ab.absxs.body_y\[4\] net869 net963 _03216_ _08264_ vssd1
+ vssd1 vccd1 vccd1 _08265_ sky130_fd_sc_hd__a221o_1
XANTENNA__12465__A game.CPU.applesa.ab.absxs.body_x\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09758__B game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13342_ _06597_ _06603_ _06654_ _06602_ net695 net476 vssd1 vssd1 vccd1 vccd1 _07216_
+ sky130_fd_sc_hd__mux4_1
X_16130_ _01750_ _01751_ _01752_ _01757_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__or4_1
X_10554_ game.CPU.applesa.ab.absxs.body_x\[29\] _04647_ _04650_ net930 vssd1 vssd1
+ vccd1 vccd1 _01164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12184__B net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_297_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_350_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_295_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ net501 _07144_ _07146_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__a21o_1
XANTENNA__13599__S0 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16061_ game.CPU.applesa.ab.check_walls.above.walls\[192\] net354 vssd1 vssd1 vccd1
+ vccd1 _02073_ sky130_fd_sc_hd__xnor2_1
X_10485_ game.CPU.applesa.ab.absxs.body_x\[87\] _04610_ _04611_ game.CPU.applesa.ab.absxs.body_x\[83\]
+ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12224_ net812 net419 vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__xnor2_1
X_15012_ net1220 net1248 game.CPU.applesa.ab.check_walls.above.walls\[40\] vssd1 vssd1
+ vccd1 vccd1 _00230_ sky130_fd_sc_hd__and3_1
XANTENNA__13912__B2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_324_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19820_ clknet_leaf_37_clk game.writer.tracker.next_frame\[415\] net1350 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[415\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18926__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12155_ net823 net388 vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17991__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16457__A3 _02413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14468__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11106_ _03346_ net405 vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__xnor2_1
X_19751_ clknet_leaf_25_clk game.writer.tracker.next_frame\[346\] net1321 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[346\] sky130_fd_sc_hd__dfrtp_1
X_16963_ _02423_ net94 _02659_ net1548 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[314\]
+ sky130_fd_sc_hd__a22o_1
X_12086_ _05970_ _05971_ _05972_ _05969_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__a211o_1
XANTENNA__13676__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18702_ clknet_leaf_31_clk _01119_ _00439_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[56\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_246_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11037_ game.CPU.applesa.ab.absxs.body_x\[65\] net412 net546 game.CPU.applesa.ab.absxs.body_x\[67\]
+ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__a2bb2o_1
X_15914_ game.CPU.applesa.ab.check_walls.above.walls\[134\] net438 vssd1 vssd1 vccd1
+ vccd1 _01926_ sky130_fd_sc_hd__nor2_1
X_19682_ clknet_leaf_34_clk game.writer.tracker.next_frame\[277\] net1338 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[277\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16400__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16894_ _02464_ net93 _02640_ net1700 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[264\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_246_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18595__Q game.CPU.applesa.ab.absxs.body_y\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18633_ clknet_leaf_11_clk _01050_ _00370_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_15845_ _03387_ net353 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11544__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15016__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18564_ clknet_leaf_13_clk _00984_ _00301_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[117\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15776_ _03254_ net351 net462 game.CPU.applesa.ab.absxs.body_x\[107\] _01787_ vssd1
+ vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a221o_1
X_12988_ game.writer.tracker.frame\[554\] game.writer.tracker.frame\[555\] net1006
+ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_335_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12359__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17515_ _02883_ _02911_ _02915_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__or3_1
X_14727_ _03505_ _08557_ vssd1 vssd1 vccd1 vccd1 _08559_ sky130_fd_sc_hd__nor2_1
XANTENNA__16917__A1 _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11939_ net748 _05587_ _05589_ net572 _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__o221a_1
X_18495_ net599 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__inv_2
XANTENNA__11454__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12651__B2 game.CPU.applesa.ab.absxs.body_y\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18327__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17446_ _02772_ _02779_ _02817_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14658_ _04356_ _08492_ vssd1 vssd1 vccd1 vccd1 _08497_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12939__C1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13609_ net223 _07482_ vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__nand2_1
X_17377_ net1119 _02806_ _02804_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12375__A game.CPU.applesa.ab.absxs.body_x\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14589_ game.CPU.clock1.counter\[13\] _08445_ _08450_ _08440_ _08442_ vssd1 vssd1
+ vccd1 vccd1 _08451_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_15_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_305_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19116_ net1182 _00156_ _00787_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[161\]
+ sky130_fd_sc_hd__dfrtp_4
X_16328_ net238 _02320_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__nor2_4
XFILLER_0_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19701__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_298_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10607__B _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_320_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19047_ net1186 _00279_ _00718_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_298_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16259_ net235 _02264_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__nand2_1
XANTENNA__14590__A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire755_A _03528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09684__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19851__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14459__A2 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19949_ clknet_leaf_38_clk game.writer.tracker.next_frame\[544\] net1334 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[544\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13667__B1 _07524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09702_ net916 game.CPU.applesa.ab.check_walls.above.walls\[57\] _03415_ net1143
+ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a22o_1
XFILLER_0_241_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13419__A0 _06649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09633_ net1084 _03282_ _03354_ net1158 _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__a221o_1
XFILLER_0_241_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout270_A game.CPU.walls.rand_wall.abduyd.next_wall\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09564_ net1106 net1267 vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__xor2_1
XFILLER_0_306_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12269__B net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11173__B net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09495_ net1133 net818 vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__nand2_1
XANTENNA__16908__B2 game.writer.tracker.frame\[273\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout156_X net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18237__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout535_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17030__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1277_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout702_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1065_X net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19381__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18949__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16687__A3 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_230_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1232_X net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13355__C1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09594__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ game.CPU.applesa.ab.collisions game.CPU.applesa.ab.check_walls.impossible
+ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10533__A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13107__C1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout440 net443 vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_306_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout957_X net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19555__RESET_B net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout451 _08425_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_6
XANTENNA__13844__A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout462 net464 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_8
Xfanout473 net474 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_8
X_13960_ net939 net783 vssd1 vssd1 vccd1 vccd1 _07834_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_144_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout484 net485 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_4
Xfanout495 net496 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_283_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout69_X net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ net490 _06784_ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__or2_1
X_13891_ _07762_ _07763_ _07764_ _07761_ vssd1 vssd1 vccd1 vccd1 _07765_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_241_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11364__A game.CPU.applesa.ab.check_walls.above.walls\[35\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15630_ game.CPU.applesa.ab.check_walls.above.walls\[184\] net354 net450 net782 _01641_
+ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__a221o_1
X_12842_ game.writer.tracker.frame\[274\] game.writer.tracker.frame\[275\] net1018
+ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15561_ _08936_ _01579_ _01578_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12633__A1 game.CPU.applesa.ab.absxs.body_x\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12773_ game.writer.tracker.frame\[86\] game.writer.tracker.frame\[87\] net1028 vssd1
+ vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__mux2_1
XANTENNA__12894__S net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13830__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12633__B2 game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17300_ net2029 net721 _02756_ _02383_ net175 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[554\]
+ sky130_fd_sc_hd__a32o_1
X_14512_ game.CPU.apple_location2\[1\] net881 net856 game.CPU.apple_location2\[7\]
+ vssd1 vssd1 vccd1 vccd1 _08386_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_25_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ net751 _05332_ _05337_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a21oi_1
X_18280_ net622 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
XANTENNA__09769__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_327_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15492_ _08404_ _01515_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__nand2_4
XANTENNA__19724__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14394__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17572__A1 _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17231_ _02544_ net78 _02738_ net1695 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[503\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14443_ net1268 net1045 vssd1 vssd1 vccd1 vccd1 _08317_ sky130_fd_sc_hd__or2_1
XANTENNA__17986__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11655_ game.CPU.applesa.ab.check_walls.above.walls\[12\] net252 _05543_ vssd1 vssd1
+ vccd1 vccd1 _05544_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_299_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12195__A game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15583__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout80 net82 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_2
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_330_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout91 _02637_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__buf_4
X_17162_ net149 _02452_ net77 _02721_ net1501 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[451\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10606_ _04174_ _04583_ _04591_ _04625_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a31o_4
X_14374_ game.CPU.applesa.ab.absxs.body_y\[119\] net946 vssd1 vssd1 vccd1 vccd1 _08248_
+ sky130_fd_sc_hd__xor2_1
X_11586_ game.CPU.applesa.ab.check_walls.above.walls\[108\] net251 vssd1 vssd1 vccd1
+ vccd1 _05475_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16127__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15002__C game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_302_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13578__X _07452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16113_ game.CPU.applesa.ab.absxs.body_y\[68\] net452 vssd1 vssd1 vccd1 vccd1 _02125_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__14138__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13325_ net211 _07198_ _07197_ net277 vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__a211o_1
XANTENNA__14138__B2 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10537_ game.CPU.applesa.ab.absxs.body_x\[45\] _04640_ _04641_ game.CPU.applesa.ab.absxs.body_x\[41\]
+ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__a22o_1
X_17093_ _02327_ net58 _02699_ net1652 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[404\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19874__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12923__A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13346__C1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16044_ game.CPU.applesa.ab.absxs.body_x\[47\] net463 net442 game.CPU.applesa.ab.absxs.body_y\[46\]
+ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a22o_1
X_13256_ game.writer.tracker.frame\[456\] game.writer.tracker.frame\[457\] net1014
+ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__mux2_1
X_10468_ net931 game.CPU.applesa.ab.absxs.body_x\[96\] _04594_ _04599_ vssd1 vssd1
+ vccd1 vccd1 _01199_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_94_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13361__A2 _06678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12207_ _05922_ _06092_ _05920_ _05921_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__or4bb_1
X_13187_ game.writer.tracker.frame\[436\] game.writer.tracker.frame\[437\] net1036
+ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__mux2_1
X_10399_ net1260 _04358_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_244_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11372__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19803_ clknet_leaf_33_clk game.writer.tracker.next_frame\[398\] net1324 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[398\] sky130_fd_sc_hd__dfrtp_1
X_12138_ game.CPU.applesa.ab.check_walls.above.walls\[71\] net297 net292 net814 _06024_
+ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__a221o_1
XANTENNA__15953__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13649__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17995_ net656 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__inv_2
XANTENNA__16401__Y _02373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_341_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19734_ clknet_leaf_19_clk game.writer.tracker.next_frame\[329\] net1317 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[329\] sky130_fd_sc_hd__dfrtp_2
X_16946_ _02390_ net87 _02654_ net1728 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[301\]
+ sky130_fd_sc_hd__a22o_1
X_12069_ game.CPU.applesa.ab.check_walls.above.walls\[124\] net551 vssd1 vssd1 vccd1
+ vccd1 _05956_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_223_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_193_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_251_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19665_ clknet_leaf_30_clk game.writer.tracker.next_frame\[260\] net1291 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[260\] sky130_fd_sc_hd__dfrtp_1
X_16877_ _02438_ net122 _02630_ game.writer.tracker.frame\[257\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[257\] sky130_fd_sc_hd__a22o_1
XFILLER_0_223_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11675__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19214__Q game.CPU.applesa.ab.apple_possible\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18616_ clknet_leaf_13_clk _01033_ _00353_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[110\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16602__A3 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10883__B1 game.CPU.applesa.ab.apple_possible\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15828_ game.CPU.applesa.ab.absxs.body_y\[19\] net433 vssd1 vssd1 vccd1 vccd1 _01840_
+ sky130_fd_sc_hd__xnor2_1
X_19596_ clknet_leaf_36_clk game.writer.tracker.next_frame\[191\] net1355 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[191\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14074__B1 game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16784__B net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12089__B net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18547_ net633 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__inv_2
X_15759_ game.CPU.applesa.ab.absxs.body_y\[23\] net433 vssd1 vssd1 vccd1 vccd1 _01771_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_47_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17012__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_255_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09679__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09280_ game.CPU.applesa.twomode.counter_normal vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__inv_2
X_18478_ net636 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_333_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_177_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17429_ _03219_ _02832_ _02835_ _02853_ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a31o_1
XANTENNA__09398__B net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_306_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10938__A1 game.CPU.applesa.ab.absxs.body_x\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10938__B2 game.CPU.applesa.ab.absxs.body_y\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_259_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13929__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10905__X _00015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout116_A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16305__A _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload50 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 clkload50/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_286_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload61 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_286_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload72 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__inv_6
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12552__B net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09556__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16024__B net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_266_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09556__B2 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10353__A game.CPU.walls.rand_wall.input2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1025_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11363__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11363__B2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11168__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15863__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ game.CPU.applesa.ab.absxs.body_x\[38\] vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout485_A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16841__A3 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16040__A game.CPU.applesa.ab.absxs.body_x\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout273_X net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16054__A1 game.CPU.applesa.ab.absxs.body_x\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_183_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16054__B2 game.CPU.applesa.ab.absxs.body_y\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09616_ net1140 game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1
+ vccd1 _03859_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_355_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18621__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19747__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09547_ net1160 game.CPU.applesa.ab.absxs.body_y\[112\] vssd1 vssd1 vccd1 vccd1 _03790_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_203_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14495__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_277_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout917_A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16357__A2 _02258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ net1108 game.CPU.applesa.ab.check_walls.above.walls\[176\] vssd1 vssd1 vccd1
+ vccd1 _03721_ sky130_fd_sc_hd__xor2_1
XFILLER_0_337_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_175_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18771__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19897__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12379__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload0 clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__inv_12
XANTENNA__09876__X _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11440_ game.CPU.applesa.ab.check_walls.above.walls\[30\] net256 vssd1 vssd1 vccd1
+ vccd1 _05329_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13040__A1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09795__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11371_ net745 _05255_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__nor2_1
XANTENNA__09795__B2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16215__A _06571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19127__CLK net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13110_ _06976_ _06982_ _06983_ net186 vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__a211o_1
X_10322_ game.CPU.randy.f1.a1.count\[11\] _04500_ net1988 vssd1 vssd1 vccd1 vccd1
+ _04502_ sky130_fd_sc_hd__a21oi_1
X_14090_ net1058 game.CPU.applesa.ab.check_walls.above.walls\[10\] vssd1 vssd1 vccd1
+ vccd1 _07964_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_308_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12462__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10534__Y _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13041_ net481 _06912_ _06914_ net282 vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_150_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10253_ net569 _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__nand2_1
XFILLER_0_277_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11078__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15773__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ net1125 _04375_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__nor2_1
Xfanout1202 game.CPU.walls.rand_wall.good_spot vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__buf_2
XFILLER_0_292_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1213 net1214 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__clkbuf_2
XANTENNA__19277__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1224 net1228 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__clkbuf_2
X_16800_ net157 _02322_ net99 net730 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__o31a_1
XFILLER_0_273_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1235 net1236 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16588__C _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1246 net1247 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__dlymetal6s2s_1
X_17780_ game.CPU.applesa.twoapples.count\[1\] _03125_ _03129_ vssd1 vssd1 vccd1 vccd1
+ _03130_ sky130_fd_sc_hd__o21ai_1
XANTENNA__16832__A3 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14992_ net1224 net1255 game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1
+ vccd1 vccd1 _00208_ sky130_fd_sc_hd__and3_1
Xfanout1257 game.CPU.walls.enable_in vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__buf_4
Xfanout1268 game.CPU.applesa.ab.absxs.body_x\[91\] vssd1 vssd1 vccd1 vccd1 net1268
+ sky130_fd_sc_hd__clkbuf_2
Xfanout270 game.CPU.walls.rand_wall.abduyd.next_wall\[0\] vssd1 vssd1 vccd1 vccd1
+ net270 sky130_fd_sc_hd__buf_4
Xfanout281 net282 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13500__C1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1279 net1280 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__clkbuf_4
X_16731_ _02561_ _02579_ net718 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__o21a_1
Xfanout292 _05861_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_4
X_13943_ net1048 _03417_ game.CPU.applesa.ab.check_walls.above.walls\[69\] net864
+ _07815_ vssd1 vssd1 vccd1 vccd1 _07817_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19450_ clknet_leaf_47_clk game.writer.tracker.next_frame\[45\] net1299 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[45\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16662_ net152 net129 _02428_ _02548_ net1659 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[124\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13874_ net1061 game.CPU.applesa.ab.check_walls.above.walls\[105\] vssd1 vssd1 vccd1
+ vccd1 _07748_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16596__A2 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17793__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13912__A1_N net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_319_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18401_ net617 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__inv_2
X_15613_ net810 net451 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__xnor2_1
X_12825_ game.writer.tracker.frame\[358\] game.writer.tracker.frame\[359\] net1001
+ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__mux2_1
X_19381_ clknet_leaf_10_clk _01387_ _00961_ vssd1 vssd1 vccd1 vccd1 game.CPU.bodymain1.main.score\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_16593_ net1819 _02505_ _02508_ net126 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[95\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13803__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18332_ net594 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15544_ net954 _01545_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09499__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12756_ game.writer.tracker.frame\[110\] game.writer.tracker.frame\[111\] net995
+ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09483__B1 game.CPU.applesa.ab.check_walls.above.walls\[178\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17545__A1 _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Left_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11541__B net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11707_ net787 net254 vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15013__B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11290__B1 _05178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18263_ net648 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__inv_2
XANTENNA__16899__A3 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15475_ _01454_ _01488_ _01485_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__a21o_1
X_12687_ _06559_ _06560_ _06558_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_56_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17214_ _02533_ net75 _02734_ net1862 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[490\]
+ sky130_fd_sc_hd__a22o_1
X_14426_ _08293_ _08294_ _08296_ vssd1 vssd1 vccd1 vccd1 _08300_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11638_ net774 _05526_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18194_ net608 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__inv_2
XANTENNA__15948__B net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17145_ net185 _02418_ net80 _02715_ net1649 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[440\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13582__A2 game.writer.tracker.frame\[376\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14357_ game.CPU.applesa.ab.absxs.body_y\[100\] net985 vssd1 vssd1 vccd1 vccd1 _08231_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_250_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11569_ _05457_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13308_ net224 _07177_ _07181_ net281 vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__a211o_1
X_17076_ net216 _02373_ net60 _02695_ net1756 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[391\]
+ sky130_fd_sc_hd__a32o_1
X_14288_ game.CPU.applesa.ab.absxs.body_x\[84\] net886 net1060 _03233_ vssd1 vssd1
+ vccd1 vccd1 _08162_ sky130_fd_sc_hd__o22a_1
XANTENNA__16520__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19209__Q game.CPU.applesa.ab.apple_possible\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16027_ _02035_ _02036_ _02037_ _02038_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__or4_1
XFILLER_0_295_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13239_ _07109_ _07110_ _07112_ _07111_ net489 net683 vssd1 vssd1 vccd1 vccd1 _07113_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_268_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Left_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16808__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__B1 game.CPU.applesa.twoapples.absxs.next_head\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17076__A3 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15683__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13717__S0 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17978_ net607 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14295__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18644__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_305_Left_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19717_ clknet_leaf_35_clk game.writer.tracker.next_frame\[312\] net1345 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[312\] sky130_fd_sc_hd__dfrtp_1
X_16929_ _02512_ net97 _02650_ game.writer.tracker.frame\[289\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[289\] sky130_fd_sc_hd__a22o_1
XFILLER_0_251_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09710__A1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09710__B2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19648_ clknet_leaf_21_clk game.writer.tracker.next_frame\[243\] net1337 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[243\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16587__A2 _02387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_179_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ net1101 _03428_ game.CPU.applesa.ab.check_walls.above.walls\[90\] net922
+ _03639_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__a221o_1
XANTENNA__18783__Q game.CPU.applesa.ab.absxs.body_x\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13931__B net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19579_ clknet_leaf_32_clk game.writer.tracker.next_frame\[174\] net1284 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[174\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18794__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15795__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_124_Left_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11291__X _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09332_ net1090 _03265_ game.CPU.applesa.ab.absxs.body_y\[82\] net902 vssd1 vssd1
+ vccd1 vccd1 _03575_ sky130_fd_sc_hd__a22o_1
XANTENNA__13270__A1 game.writer.tracker.frame\[497\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09474__B1 game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12547__B net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11762__A1_N net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16019__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09202__A game.CPU.applesa.ab.check_walls.above.walls\[135\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11281__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ game.CPU.randy.counter1.count1\[4\] vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout233_A _04701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11820__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_350_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_314_Left_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09194_ net796 vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_306_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09856__B game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16035__A game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1142_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout119_X net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12282__B net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09529__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19119__Q game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_133_Left_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09529__B2 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12850__X _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18250__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12533__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18958__Q game.CPU.applesa.ab.check_walls.above.walls\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_328_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 game.writer.control.button5.Q\[1\] vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_323_Left_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold23 game.CPU.right_button.eD1.Q1 vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13089__A1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_227_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_328_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold34 game.CPU.walls.abc.number\[6\] vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14286__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ game.CPU.applesa.ab.absxs.body_x\[102\] vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_303_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold45 game.CPU.applesa.ab.y_final\[0\] vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_270_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold56 game.CPU.applesa.ab.x_final\[0\] vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_279_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold67 game.writer.tracker.frame\[140\] vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold78 game.CPU.applesa.apple_location2_n\[5\] vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 game.writer.tracker.frame\[47\] vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17224__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09701__A1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10940_ _04820_ _04829_ _04826_ _04828_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__or4b_1
XANTENNA__09701__B2 net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18693__Q game.CPU.applesa.ab.absxs.body_x\[35\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_357_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871_ _04767_ _04773_ game.CPU.randy.counter1.count\[18\] _03495_ vssd1 vssd1 vccd1
+ vccd1 _04774_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_280_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12610_ _06251_ _06258_ _06349_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_344_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13590_ game.writer.tracker.frame\[345\] game.writer.tracker.frame\[347\] game.writer.tracker.frame\[348\]
+ game.writer.tracker.frame\[346\] net975 net1018 vssd1 vssd1 vccd1 vccd1 _07464_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_195_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_356_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09112__A net1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11361__B net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_332_Left_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12541_ game.CPU.applesa.ab.absxs.body_x\[42\] net371 net360 game.CPU.applesa.ab.absxs.body_y\[40\]
+ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__a22o_1
XANTENNA__10258__A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_314_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_352_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15260_ _08817_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
XFILLER_0_289_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12472_ _06343_ _06344_ _06345_ _06348_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_152_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08951__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16750__A2 _02391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14211_ game.CPU.applesa.ab.absxs.body_y\[92\] net983 vssd1 vssd1 vccd1 vccd1 _08085_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__13564__A2 _07429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11423_ net796 net259 _05311_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a21oi_1
X_15191_ _04587_ _04628_ _08755_ vssd1 vssd1 vccd1 vccd1 _08763_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_229_Right_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_340_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_9 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14142_ _07939_ _07940_ _07949_ _07983_ vssd1 vssd1 vccd1 vccd1 _08016_ sky130_fd_sc_hd__a31o_1
X_11354_ net563 _05236_ _05242_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19029__Q game.CPU.applesa.ab.check_walls.above.walls\[74\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10305_ game.CPU.randy.f1.a1.count\[2\] game.CPU.randy.f1.a1.count\[1\] game.CPU.randy.f1.a1.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__and3_1
X_14073_ net888 game.CPU.applesa.ab.check_walls.above.walls\[0\] _03379_ net985 vssd1
+ vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__o22a_1
X_18950_ clknet_leaf_67_clk net1400 _00621_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11285_ _05062_ _05064_ _05069_ _05071_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__or4_1
XANTENNA__16232__X _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11327__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18667__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16599__B _02512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13024_ _06861_ _06880_ net697 vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__mux2_1
X_10236_ _04363_ _04371_ _04365_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__a21o_1
XANTENNA__09782__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17901_ net639 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__inv_2
XANTENNA__19912__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18881_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[11\] _00576_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_265_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_238_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1010 net1011 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__clkbuf_4
Xfanout1021 net1022 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_4
X_17832_ game.writer.updater.commands.count\[5\] _03158_ _03150_ vssd1 vssd1 vccd1
+ vccd1 _03162_ sky130_fd_sc_hd__o21ai_1
Xfanout1032 net1033 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_4
X_10167_ _04359_ net1078 _04357_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__or3b_1
XFILLER_0_238_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__buf_4
XFILLER_0_206_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1054 game.CPU.applesa.x\[2\] vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_163_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1065 net1066 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_4
Xfanout1076 net1077 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11536__B net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17763_ game.CPU.applesa.twoapples.count_luck\[4\] _03116_ vssd1 vssd1 vccd1 vccd1
+ _03118_ sky130_fd_sc_hd__or2_1
X_14975_ net1225 net1253 game.CPU.applesa.ab.check_walls.above.walls\[3\] vssd1 vssd1
+ vccd1 vccd1 _00110_ sky130_fd_sc_hd__and3_1
Xfanout1087 net1088 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_4
X_10098_ game.CPU.applesa.twoapples.count_luck\[5\] game.CPU.applesa.twoapples.count_luck\[4\]
+ game.CPU.applesa.twoapples.count_luck\[1\] _04303_ vssd1 vssd1 vccd1 vccd1 _04306_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__15008__B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1098 net1099 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__clkbuf_8
X_16714_ _02336_ net100 net736 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__o21a_1
X_19502_ clknet_leaf_27_clk game.writer.tracker.next_frame\[97\] net1309 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[97\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_254_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13926_ net941 game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1 vccd1
+ vccd1 _07800_ sky130_fd_sc_hd__xor2_1
XFILLER_0_261_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14029__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17694_ _03062_ _03073_ _03074_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__nor3_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19433_ clknet_leaf_41_clk game.writer.tracker.next_frame\[28\] net1352 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_254_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16645_ net1785 _02540_ _02541_ net126 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[114\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17230__A3 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13857_ game.writer.tracker.frame\[545\] game.writer.tracker.frame\[547\] game.writer.tracker.frame\[548\]
+ game.writer.tracker.frame\[546\] net971 net1006 vssd1 vssd1 vccd1 vccd1 _07731_
+ sky130_fd_sc_hd__mux4_1
X_12808_ _06678_ _06679_ _06681_ _06680_ net478 net678 vssd1 vssd1 vccd1 vccd1 _06682_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19364_ clknet_leaf_69_clk _01370_ _00945_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_16576_ _02356_ _02376_ vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__nor2_4
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13788_ game.writer.tracker.frame\[393\] game.writer.tracker.frame\[395\] game.writer.tracker.frame\[396\]
+ game.writer.tracker.frame\[394\] net977 net1020 vssd1 vssd1 vccd1 vccd1 _07662_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_44_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17518__B2 net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_252_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18315_ net620 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__inv_2
XANTENNA__09022__A game.CPU.applesa.ab.absxs.body_x\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15527_ _01474_ _01548_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12739_ net488 _06612_ net686 vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__a21o_1
XANTENNA__15959__A game.CPU.applesa.ab.check_walls.above.walls\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_19295_ clknet_leaf_68_clk _01339_ _00914_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.logic_enable
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18335__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09957__A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18246_ net644 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
X_15458_ _01456_ _01483_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15678__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14201__B1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12654__Y _06531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19442__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11015__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14409_ game.CPU.applesa.ab.absxs.body_x\[44\] net890 net952 _03309_ vssd1 vssd1
+ vccd1 vccd1 _08283_ sky130_fd_sc_hd__a22o_1
XANTENNA__10455__X _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18177_ net609 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__inv_2
XANTENNA__09676__B game.CPU.applesa.ab.absxs.body_y\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15389_ _08903_ _08920_ vssd1 vssd1 vccd1 vccd1 _08931_ sky130_fd_sc_hd__or2_2
XANTENNA__12383__A game.CPU.applesa.ab.absxs.body_y\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold504 game.writer.tracker.frame\[83\] vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
X_17128_ game.writer.tracker.frame\[428\] _02710_ vssd1 vssd1 vccd1 vccd1 _02711_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_80_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15800__A2_N net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold515 game.CPU.applesa.apple_location2_n\[2\] vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_279_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold526 game.writer.tracker.frame\[269\] vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold537 game.writer.tracker.frame\[464\] vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 game.CPU.randy.f1.a1.count\[11\] vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
X_17059_ _02429_ net83 _02688_ net1620 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[381\]
+ sky130_fd_sc_hd__a22o_1
Xhold559 game.writer.tracker.frame\[325\] vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09950_ _04175_ _04177_ _04183_ vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__o21a_1
XFILLER_0_311_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10107__S _04311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19592__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_263_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09692__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09881_ _03836_ _03839_ _03847_ _03774_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__o31a_1
XANTENNA__13926__B game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16302__B net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload18_A clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_295_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14268__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14103__A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout183_A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13942__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_352_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17221__A3 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15768__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout350_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19402__Q game.CPU.applesa.x\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1092_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout448_A _08427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_274_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_314_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09447__B1 game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16980__A2 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11254__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09315_ net1086 game.CPU.applesa.ab.absxs.body_x\[67\] vssd1 vssd1 vccd1 vccd1 _03558_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__11181__B net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_216_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout615_A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18245__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09867__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09246_ game.CPU.applesa.ab.good_spot vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16193__B1 _02196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_330_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09177_ net808 vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12293__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1145_X net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11557__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Left_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_322_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19935__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout984_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput13 net13 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
Xoutput35 net35 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_285_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XANTENNA_fanout96_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11070_ game.CPU.applesa.ab.absxs.body_x\[27\] net546 net541 game.CPU.applesa.ab.absxs.body_y\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_227_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15891__X _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ net1125 _04226_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__nor2_1
XANTENNA__14013__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09107__A game.CPU.applesa.ab.absxs.body_y\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__B net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12904__S1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14760_ game.CPU.randy.counter1.count\[15\] net265 _03499_ vssd1 vssd1 vccd1 vccd1
+ _08581_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13482__A1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ _05855_ _05856_ net293 net789 _05857_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a221o_1
XFILLER_0_291_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13711_ _07583_ _07584_ net478 vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_2_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923_ net1166 _04362_ _04813_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_316_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _04351_ net752 vssd1 vssd1 vccd1 vccd1 _08530_ sky130_fd_sc_hd__nor2_1
XANTENNA__12468__A game.CPU.applesa.ab.absxs.body_y\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16420__A1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_296_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16430_ net115 net164 net67 _02388_ net1474 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[47\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13642_ _07514_ _07515_ net499 vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10854_ _04756_ _04755_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_238_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14431__B1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16971__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16882__B net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12187__B net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11091__B net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16361_ net181 _02241_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__nand2_4
XANTENNA__11245__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13573_ game.writer.tracker.frame\[357\] game.writer.tracker.frame\[359\] game.writer.tracker.frame\[360\]
+ game.writer.tracker.frame\[358\] net968 net1001 vssd1 vssd1 vccd1 vccd1 _07447_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ game.CPU.applesa.ab.absxs.body_y\[51\] _04630_ vssd1 vssd1 vccd1 vccd1 _04724_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11796__A1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18100_ net614 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__inv_2
X_15312_ _08858_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09777__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19080_ net1179 _00116_ _00751_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12524_ game.CPU.applesa.ab.absxs.body_y\[71\] net365 vssd1 vssd1 vccd1 vccd1 _06401_
+ sky130_fd_sc_hd__xnor2_1
X_16292_ net1909 net720 _02292_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[10\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__16723__A2 _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15526__A3 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_240_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18031_ net590 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15243_ game.CPU.kyle.L1.cnt_500hz\[5\] game.CPU.kyle.L1.cnt_500hz\[4\] _08802_ vssd1
+ vssd1 vccd1 vccd1 _08804_ sky130_fd_sc_hd__and3_1
XANTENNA__09496__B net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12455_ _03271_ game.CPU.applesa.twoapples.absxs.next_head\[3\] net526 game.CPU.applesa.ab.absxs.body_y\[49\]
+ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__a221o_1
XFILLER_0_297_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_229_Left_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11548__B2 game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11406_ _05280_ _05281_ _05293_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15174_ _08749_ vssd1 vssd1 vccd1 vccd1 _08750_ sky130_fd_sc_hd__inv_2
XANTENNA__15010__C net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12386_ game.CPU.applesa.ab.absxs.body_x\[24\] net385 vssd1 vssd1 vccd1 vccd1 _06263_
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_327_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14125_ net889 game.CPU.applesa.ab.check_walls.above.walls\[24\] game.CPU.applesa.ab.check_walls.above.walls\[25\]
+ net885 vssd1 vssd1 vccd1 vccd1 _07999_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11337_ game.CPU.applesa.ab.check_walls.above.walls\[82\] net767 vssd1 vssd1 vccd1
+ vccd1 _05226_ sky130_fd_sc_hd__xor2_2
XANTENNA__12931__A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19982_ clknet_leaf_44_clk _01406_ net1298 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_265_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14498__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_238_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10771__A2 _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14056_ net938 net789 vssd1 vssd1 vccd1 vccd1 _07930_ sky130_fd_sc_hd__xor2_1
X_18933_ clknet_leaf_5_clk net1388 _00617_ vssd1 vssd1 vccd1 vccd1 game.CPU.start_pause_button1.eD1.D
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18598__Q game.CPU.applesa.ab.absxs.body_y\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11268_ _04858_ _04861_ _05156_ _05157_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__or4_1
XANTENNA__13170__B1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13238__S net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13007_ game.writer.tracker.frame\[556\] game.writer.tracker.frame\[557\] net1006
+ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__mux2_1
X_10219_ _04408_ _04411_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15019__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18864_ clknet_leaf_0_clk _01255_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11199_ game.CPU.applesa.ab.absxs.body_x\[23\] net544 net538 game.CPU.applesa.ab.absxs.body_y\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__a22o_1
X_17815_ _03149_ game.writer.updater.commands.count\[0\] net182 vssd1 vssd1 vccd1
+ vccd1 _01409_ sky130_fd_sc_hd__mux2_1
XANTENNA__15961__B net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15998__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18795_ clknet_leaf_4_clk _01210_ _00532_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_238_Left_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17746_ game.CPU.applesa.ab.good_collision net851 _03103_ game.CPU.applesa.ab.start_enable
+ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__o211a_1
X_14958_ _08660_ _08664_ _08734_ _08705_ vssd1 vssd1 vccd1 vccd1 _08735_ sky130_fd_sc_hd__o31a_1
XFILLER_0_89_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13473__A1 _07096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_338_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13909_ net881 game.CPU.applesa.ab.check_walls.above.walls\[121\] _03446_ net948
+ _07782_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17203__A3 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17677_ _03062_ _03063_ _03064_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__nor3_1
XFILLER_0_159_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14889_ net1090 _08419_ vssd1 vssd1 vccd1 vccd1 _08666_ sky130_fd_sc_hd__nor2_1
XANTENNA__19808__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16411__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16628_ _02381_ _02520_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__nor2_2
X_19416_ clknet_leaf_48_clk game.writer.tracker.next_frame\[11\] net1296 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14422__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19839__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16559_ net151 _02486_ vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__and2_1
X_19347_ clknet_leaf_72_clk game.CPU.applesa.twoapples.good_spot_next vssd1 vssd1
+ vccd1 vccd1 game.CPU.applesa.twoapples.good_spot sky130_fd_sc_hd__dfxtp_1
XFILLER_0_335_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09100_ game.CPU.applesa.ab.absxs.body_y\[26\] vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__inv_2
XANTENNA__10329__C net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12984__B1 _06639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19278_ clknet_leaf_7_clk _00048_ _00908_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__19958__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16714__A2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09031_ game.CPU.applesa.ab.absxs.body_x\[25\] vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18229_ net665 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_349_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold301 game.writer.tracker.frame\[483\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_211_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold312 game.writer.tracker.frame\[360\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 game.writer.tracker.frame\[275\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_269_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold334 game.writer.tracker.frame\[112\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16478__B2 _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18982__CLK net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 game.writer.tracker.frame\[108\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16313__A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold356 game.writer.tracker.frame\[228\] vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14489__B1 _08062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold367 game.writer.tracker.frame\[39\] vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10762__A2 _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold378 game.writer.tracker.frame\[208\] vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 game.writer.tracker.frame\[455\] vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net1109 net847 _04171_ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_6_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout803 game.CPU.applesa.ab.check_walls.above.walls\[102\] vssd1 vssd1 vccd1 vccd1
+ net803 sky130_fd_sc_hd__buf_2
Xfanout814 game.CPU.applesa.ab.check_walls.above.walls\[70\] vssd1 vssd1 vccd1 vccd1
+ net814 sky130_fd_sc_hd__buf_4
XFILLER_0_68_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_284_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout825 game.CPU.applesa.ab.check_walls.above.walls\[31\] vssd1 vssd1 vccd1 vccd1
+ net825 sky130_fd_sc_hd__buf_4
XFILLER_0_309_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout398_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20053_ net1371 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
Xfanout836 net840 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_2
XANTENNA__09904__B2 net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09864_ net900 game.CPU.applesa.ab.absxs.body_y\[45\] game.CPU.applesa.ab.absxs.body_y\[44\]
+ net894 _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__a221o_1
Xfanout847 net849 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__buf_2
XFILLER_0_244_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout858 net859 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__clkbuf_4
XANTENNA__19338__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1105_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10514__A2 _03527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout869 _03374_ vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__buf_4
XFILLER_0_99_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11176__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15871__B net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09795_ net1084 _03274_ game.CPU.applesa.ab.absxs.body_x\[42\] net922 _04037_ vssd1
+ vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_300_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout186_X net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16650__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_240_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_222_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19488__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19132__Q game.CPU.applesa.ab.check_walls.above.walls\[177\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12288__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1095_X net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14413__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13767__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11778__B2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10570_ net1123 game.CPU.bodymain1.main.score\[0\] _04656_ _04594_ vssd1 vssd1 vccd1
+ vccd1 _04657_ sky130_fd_sc_hd__o31a_2
XANTENNA__09597__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16705__A2 _02486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_311_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1 vssd1 vccd1 vccd1
+ _03478_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_233_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09884__X _04127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12240_ game.CPU.applesa.ab.check_walls.above.walls\[151\] net422 vssd1 vssd1 vccd1
+ vccd1 _06126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14192__A2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout987_X net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16469__B2 _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ _06055_ _06056_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__or3_1
XFILLER_0_247_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17130__A2 _02387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout99_X net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10753__A2 _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11122_ game.CPU.applesa.ab.absxs.body_y\[18\] net401 vssd1 vssd1 vccd1 vccd1 _05012_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_219_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11053_ _03255_ net324 vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__xnor2_1
X_15930_ game.CPU.applesa.ab.check_walls.above.walls\[124\] net449 vssd1 vssd1 vccd1
+ vccd1 _01942_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10271__A game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11702__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10505__A2 _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10004_ net1165 game.CPU.applesa.out_random_2\[0\] vssd1 vssd1 vccd1 vccd1 _04212_
+ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_322_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11086__B net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15861_ game.CPU.applesa.ab.absxs.body_x\[113\] net473 vssd1 vssd1 vccd1 vccd1 _01873_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12897__S net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18705__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17600_ game.CPU.kyle.L1.cnt_20ms\[4\] _03002_ game.CPU.kyle.L1.cnt_20ms\[5\] vssd1
+ vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08947__Y _03197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16641__A1 game.writer.tracker.frame\[113\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14812_ game.CPU.randy.counter1.count\[12\] _08619_ net138 vssd1 vssd1 vccd1 vccd1
+ _08622_ sky130_fd_sc_hd__o21ai_1
XANTENNA__16641__B2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18580_ clknet_leaf_53_clk _01000_ _00317_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[41\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13455__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15792_ _01797_ _01798_ _01802_ _01803_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__a211o_1
XANTENNA__14397__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17531_ net1259 _02875_ _02956_ _02957_ _02958_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11814__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14743_ game.CPU.randy.counter1.count1\[13\] _08567_ vssd1 vssd1 vccd1 vccd1 _08570_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_203_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11955_ _05834_ _05839_ _05842_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__and3_1
XANTENNA__17197__A2 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19042__Q game.CPU.applesa.ab.check_walls.above.walls\[87\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12198__A game.CPU.applesa.ab.check_walls.above.walls\[53\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10906_ game.CPU.modea.Qa\[0\] game.CPU.applesa.enable_in _04735_ vssd1 vssd1 vccd1
+ vccd1 _00009_ sky130_fd_sc_hd__mux2_1
X_17462_ _02785_ _02791_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__nand2_1
XANTENNA__13207__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14674_ game.CPU.randy.counter1.count1\[4\] _04347_ _08511_ _08512_ vssd1 vssd1 vccd1
+ vccd1 _08513_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_28_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15005__C game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11886_ net574 _05351_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_357_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_345_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16413_ net203 _02381_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__nor2_4
XFILLER_0_184_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19201_ clknet_leaf_67_clk _01310_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13625_ game.writer.tracker.frame\[305\] game.writer.tracker.frame\[307\] game.writer.tracker.frame\[308\]
+ game.writer.tracker.frame\[306\] net978 net1036 vssd1 vssd1 vccd1 vccd1 _07499_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__19932__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13758__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17393_ game.CPU.clock1.game_state\[0\] _02821_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10837_ game.CPU.randy.counter1.count\[17\] _03496_ vssd1 vssd1 vccd1 vccd1 _04740_
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19132_ net1183 _00173_ _00803_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[177\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_158_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16344_ net136 _02258_ net69 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_333_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13556_ game.writer.tracker.frame\[101\] net834 net672 game.writer.tracker.frame\[104\]
+ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__o22a_1
X_10768_ game.CPU.applesa.ab.absxs.body_y\[80\] _04673_ _04674_ game.CPU.applesa.ab.absxs.body_y\[76\]
+ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__a22o_1
XANTENNA__12430__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_281_Right_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_171_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16117__B net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19063_ net1186 _00097_ _00734_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[108\]
+ sky130_fd_sc_hd__dfrtp_4
X_12507_ game.CPU.applesa.ab.absxs.body_y\[73\] net526 vssd1 vssd1 vccd1 vccd1 _06384_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_298_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16275_ _06573_ net245 _02231_ _02279_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__or4b_4
XFILLER_0_325_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13487_ net678 _07141_ _07360_ net220 vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_11_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10446__A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10699_ game.CPU.applesa.ab.absxs.body_y\[79\] _04623_ _04624_ game.CPU.applesa.ab.absxs.body_y\[75\]
+ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18014_ net639 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__inv_2
XFILLER_0_301_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15226_ game.CPU.applesa.normal1.number\[1\] _08785_ net758 vssd1 vssd1 vccd1 vccd1
+ _08791_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_313_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12438_ game.CPU.applesa.ab.absxs.body_x\[107\] net530 net520 game.CPU.applesa.ab.absxs.body_y\[106\]
+ _06314_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__o221a_1
XANTENNA__14183__A2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15956__B net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_298_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15157_ net1213 net1239 game.CPU.applesa.ab.check_walls.above.walls\[185\] vssd1
+ vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12369_ _03225_ net377 vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17121__A2 _02693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_238_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14108_ _07977_ _07978_ _07979_ _07980_ vssd1 vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19965_ clknet_leaf_43_clk game.writer.tracker.next_frame\[560\] net1327 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[560\] sky130_fd_sc_hd__dfrtp_1
X_15088_ net1211 net1237 net799 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_266_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16880__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_285_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14039_ _07909_ _07910_ _07911_ _07912_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__and4bb_1
X_18916_ clknet_leaf_5_clk net5 _00600_ vssd1 vssd1 vccd1 vccd1 game.CPU.up_button.sync1.Q
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_246_Left_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_169_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19896_ clknet_leaf_14_clk game.writer.tracker.next_frame\[491\] net1283 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[491\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09898__B1 _04139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15691__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18847_ clknet_leaf_0_clk _01238_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__19630__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16632__A1 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09580_ _03821_ _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__nand2_1
X_18778_ clknet_leaf_63_clk _01195_ _00515_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[92\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17899__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17729_ game.CPU.applesa.ab.count_luck\[5\] _03093_ net1457 vssd1 vssd1 vccd1 vccd1
+ _03096_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_19_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17188__A2 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14100__B game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_258_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19780__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16935__A2 _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10680__A1 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_271_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_255_Left_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16308__A _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout146_A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_351_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12421__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12555__B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10432__A1 _04563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19010__CLK net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1055_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09014_ game.CPU.applesa.ab.absxs.body_x\[89\] vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__inv_2
XANTENNA__14174__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15866__B net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13382__B1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold120 game.writer.tracker.frame\[410\] vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 game.writer.tracker.frame\[271\] vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10643__X _04690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold142 game.writer.tracker.frame\[346\] vssd1 vssd1 vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17112__A2 _02693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1222_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold153 game.writer.tracker.frame\[214\] vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_269_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19160__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 game.writer.tracker.frame\[122\] vssd1 vssd1 vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_282_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold175 game.writer.tracker.frame\[295\] vssd1 vssd1 vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 game.writer.tracker.frame\[311\] vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_264_Left_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold197 game.writer.tracker.frame\[474\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18728__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19127__Q game.CPU.applesa.ab.check_walls.above.walls\[172\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout600 net625 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_229_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout611 net612 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__buf_4
XANTENNA__16871__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout622 net623 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__buf_4
X_09916_ net1079 net847 vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_224_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18555__RESET_B net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout633 net651 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_2
Xfanout644 net646 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_298_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_clk_X clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_X net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout655 net658 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_2
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_4
X_20036_ net1384 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
Xfanout677 _06600_ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__clkbuf_4
XANTENNA__18966__Q game.CPU.applesa.ab.check_walls.above.walls\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09847_ net1155 game.CPU.applesa.ab.absxs.body_y\[28\] vssd1 vssd1 vccd1 vccd1 _04090_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_336_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout688 net691 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_2
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 net707 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout947_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09778_ net1138 game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1 vccd1
+ vccd1 _04021_ sky130_fd_sc_hd__xor2_1
XANTENNA__18878__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_358_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout59_A net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11634__B net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15106__B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15631__A2_N net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11740_ _04441_ _05524_ _05523_ net572 vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09879__X _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_327_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16926__A2 _02643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_273_Left_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12660__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_293_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11671_ net794 net254 _05559_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_235_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ net698 _06888_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__or2_1
XFILLER_0_181_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10622_ game.CPU.applesa.ab.absxs.body_x\[67\] _04679_ _04680_ game.CPU.applesa.ab.absxs.body_x\[63\]
+ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__a22o_1
XANTENNA__16139__B1 _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14390_ game.CPU.applesa.ab.absxs.body_x\[6\] net878 net873 game.CPU.applesa.ab.absxs.body_x\[7\]
+ vssd1 vssd1 vccd1 vccd1 _08264_ sky130_fd_sc_hd__a22o_1
XANTENNA__12412__A2 net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12465__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09120__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13341_ net202 _07210_ _07214_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__a21o_1
XFILLER_0_335_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10553_ _03280_ _04647_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__nor2_1
XANTENNA__16505__X _02450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16060_ game.CPU.applesa.ab.check_walls.above.walls\[195\] net458 vssd1 vssd1 vccd1
+ vccd1 _02072_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_297_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19503__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13272_ net478 _07145_ net681 vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__a21o_1
XANTENNA__13599__S1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10484_ net1078 _04610_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__nor2_2
XFILLER_0_267_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13373__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12176__B2 game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15011_ net1215 net1241 game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1
+ vccd1 vccd1 _00229_ sky130_fd_sc_hd__and3_1
XFILLER_0_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12223_ game.CPU.applesa.ab.check_walls.above.walls\[77\] net549 vssd1 vssd1 vccd1
+ vccd1 _06109_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_282_Left_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17103__A2 _02341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_295_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12154_ game.CPU.applesa.ab.check_walls.above.walls\[134\] net288 vssd1 vssd1 vccd1
+ vccd1 _06041_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19037__Q game.CPU.applesa.ab.check_walls.above.walls\[82\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19653__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ game.CPU.applesa.ab.absxs.body_x\[35\] net408 vssd1 vssd1 vccd1 vccd1 _04995_
+ sky130_fd_sc_hd__or2_1
X_19750_ clknet_leaf_24_clk game.writer.tracker.next_frame\[345\] net1338 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[345\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_275_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16962_ _02422_ net94 _02659_ net1734 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[313\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_235_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12085_ game.CPU.applesa.ab.check_walls.above.walls\[21\] net388 vssd1 vssd1 vccd1
+ vccd1 _05972_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09790__A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18701_ clknet_leaf_60_clk _01118_ _00438_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[51\]
+ sky130_fd_sc_hd__dfrtp_4
X_11036_ _03268_ net407 net540 game.CPU.applesa.ab.absxs.body_y\[66\] vssd1 vssd1
+ vccd1 vccd1 _04926_ sky130_fd_sc_hd__a22o_1
X_15913_ _03450_ net332 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__nor2_1
X_19681_ clknet_leaf_34_clk game.writer.tracker.next_frame\[276\] net1338 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[276\] sky130_fd_sc_hd__dfrtp_1
X_16893_ net223 _02238_ _02271_ _02529_ net713 vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__o41a_1
XFILLER_0_235_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16400__B net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11825__A game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18632_ clknet_leaf_11_clk _01049_ _00369_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_15844_ game.CPU.applesa.ab.check_walls.above.walls\[23\] net434 vssd1 vssd1 vccd1
+ vccd1 _01856_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_250_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_350_Right_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15775_ _03255_ net272 net473 game.CPU.applesa.ab.absxs.body_x\[105\] vssd1 vssd1
+ vccd1 vccd1 _01787_ sky130_fd_sc_hd__a22o_1
X_18563_ clknet_leaf_13_clk _00983_ _00300_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[116\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__15016__B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_291_Left_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12987_ game.writer.tracker.frame\[546\] game.writer.tracker.frame\[547\] net1006
+ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_335_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09789__X _04032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ net1119 _04638_ _02918_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__o21ai_1
X_14726_ net54 _08557_ _08558_ vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__and3_1
X_11938_ _05585_ _05586_ _05824_ _05825_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__and4_1
X_18494_ net618 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12651__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17445_ net1258 _02873_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14657_ game.CPU.randy.counter1.count1\[17\] _08492_ _08494_ game.CPU.randy.counter1.count1\[16\]
+ _08495_ vssd1 vssd1 vccd1 vccd1 _08496_ sky130_fd_sc_hd__a221o_1
X_11869_ _04441_ _05398_ _05401_ _05755_ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__o2111a_1
X_13608_ _07480_ _07481_ net503 vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17376_ _02803_ _02805_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14588_ game.CPU.clock1.counter\[13\] _08449_ _08447_ net1275 vssd1 vssd1 vccd1 vccd1
+ _08450_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12375__B net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_333_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16327_ _06573_ net141 _02246_ net236 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__or4_2
X_19115_ net1182 _00155_ _00786_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[160\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13539_ game.writer.tracker.frame\[118\] net843 net837 game.writer.tracker.frame\[117\]
+ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__o22a_1
XFILLER_0_200_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19183__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19046_ net1191 _00278_ _00717_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[91\]
+ sky130_fd_sc_hd__dfrtp_4
X_16258_ _06571_ _06573_ _01516_ _02263_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__a31o_1
XANTENNA__15686__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15209_ net758 _08773_ _08774_ _08775_ _08776_ vssd1 vssd1 vccd1 vccd1 _08777_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_346_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09684__B net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16189_ game.CPU.applesa.ab.absxs.body_x\[71\] net462 net446 game.CPU.applesa.ab.absxs.body_y\[69\]
+ _01634_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a221o_1
XANTENNA__10717__A2 _04609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11914__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_287_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_254_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19948_ clknet_leaf_38_clk game.writer.tracker.next_frame\[543\] net1334 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[543\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10115__S _04311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16150__X _02162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13667__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ net1113 _03410_ _03411_ net1103 _03942_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__a221o_1
XANTENNA__18786__Q game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19879_ clknet_leaf_25_clk game.writer.tracker.next_frame\[474\] net1319 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[474\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10910__Y _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17406__B net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ net926 game.CPU.applesa.ab.absxs.body_x\[19\] game.CPU.applesa.ab.absxs.body_x\[17\]
+ net916 vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__a22o_1
XANTENNA__14111__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09205__A game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09563_ _03801_ _03803_ _03805_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__or3_1
X_09494_ _03734_ _03735_ _03736_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__or3_2
XANTENNA__12642__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17030__A1 _02370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__B game.CPU.applesa.ab.absxs.body_x\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout430_A net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_42_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16038__A game.CPU.applesa.ab.absxs.body_x\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_92_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout149_X net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19526__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_322_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15592__B2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12285__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18253__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1058_X net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_230_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_320_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout897_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19676__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09594__B game.CPU.applesa.ab.absxs.body_x\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_277_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11905__A1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_245_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10533__B _04639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16844__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout430 net431 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_4
Xfanout441 net443 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_4
Xfanout452 net454 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_8
Xfanout463 net464 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_2
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout474 net475 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_144_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout485 net486 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_2
X_12910_ _06658_ _06661_ net682 vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__mux2_1
Xfanout496 net499 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
X_20019_ net1277 vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_232_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13890_ net1071 _03431_ _03435_ net940 _07756_ vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_241_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12841_ game.writer.tracker.frame\[276\] game.writer.tracker.frame\[277\] net1018
+ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__mux2_1
XANTENNA__11364__B net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15560_ _01457_ _01458_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__or2_1
X_12772_ game.writer.tracker.frame\[82\] game.writer.tracker.frame\[83\] net1028 vssd1
+ vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12633__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17021__A1 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14511_ game.CPU.apple_location2\[4\] net983 vssd1 vssd1 vccd1 vccd1 _08385_ sky130_fd_sc_hd__xor2_1
X_11723_ net575 _05338_ _05332_ net749 vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_355_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15491_ _08027_ _01513_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_25_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09769__B net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12476__A game.CPU.applesa.ab.absxs.body_y\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17230_ _02415_ _02608_ net121 _02738_ net1502 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[502\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__11380__A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14442_ net1268 net1045 vssd1 vssd1 vccd1 vccd1 _08316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_355_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14386__A2 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11654_ _05537_ _05539_ _05541_ _05542_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__or4_1
XANTENNA__10267__Y _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15583__B2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout70 _02259_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12195__B net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout81 net82 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_330_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17161_ _02450_ net77 _02721_ net1792 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[450\]
+ sky130_fd_sc_hd__a22o_1
Xfanout92 net93 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__buf_2
X_10605_ game.CPU.applesa.ab.absxs.body_x\[88\] _04590_ net329 game.CPU.applesa.ab.absxs.body_x\[84\]
+ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__a22o_1
XANTENNA__15787__A game.CPU.applesa.ab.absxs.body_x\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14373_ _03288_ net1074 net1056 _03286_ _08246_ vssd1 vssd1 vccd1 vccd1 _08247_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11585_ net801 net255 vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16112_ _03277_ net270 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__xnor2_1
X_13324_ _06705_ _06707_ _06714_ _06706_ net701 net490 vssd1 vssd1 vccd1 vccd1 _07198_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09785__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17092_ net187 _02486_ net80 _02699_ net1581 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[403\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_107_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10536_ game.CPU.applesa.ab.absxs.body_x\[46\] _04640_ _04641_ game.CPU.applesa.ab.absxs.body_x\[42\]
+ vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16043_ _03310_ net338 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_310_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13255_ net277 _07121_ _07128_ net241 vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_295_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10467_ game.CPU.applesa.ab.absxs.body_x\[100\] _04595_ vssd1 vssd1 vccd1 vccd1 _04599_
+ sky130_fd_sc_hd__and2_1
XANTENNA__13897__A1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17088__A1 _02477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12206_ game.CPU.applesa.ab.check_walls.above.walls\[141\] net547 vssd1 vssd1 vccd1
+ vccd1 _06092_ sky130_fd_sc_hd__xnor2_1
X_13186_ game.writer.tracker.frame\[440\] game.writer.tracker.frame\[441\] net1038
+ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10398_ net1260 _04341_ _04548_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__o21a_1
X_19802_ clknet_leaf_33_clk game.writer.tracker.next_frame\[397\] net1324 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[397\] sky130_fd_sc_hd__dfrtp_1
X_12137_ game.CPU.applesa.ab.check_walls.above.walls\[71\] net297 net291 net814 vssd1
+ vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__o22ai_1
XANTENNA__13649__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17994_ net656 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__inv_2
XANTENNA__10580__B1 _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_179_Left_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_166_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19733_ clknet_leaf_19_clk game.writer.tracker.next_frame\[328\] net1317 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[328\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_341_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16945_ net163 net53 net87 _02655_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[300\]
+ sky130_fd_sc_hd__a31o_1
X_12068_ _05551_ _05552_ _05553_ _05554_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__or4bb_1
X_11019_ _03263_ net414 vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__nand2_1
X_19664_ clknet_leaf_30_clk game.writer.tracker.next_frame\[259\] net1291 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[259\] sky130_fd_sc_hd__dfrtp_1
X_16876_ _02553_ net107 _02630_ net1915 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[256\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10332__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17260__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_273_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18615_ clknet_leaf_13_clk _01032_ _00352_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[109\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10883__A1 game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15827_ _03283_ net352 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__xnor2_1
X_19595_ clknet_leaf_36_clk game.writer.tracker.next_frame\[190\] net1355 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[190\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14074__A1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14074__B2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_248_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18546_ net628 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__inv_2
X_15758_ _03250_ net352 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19549__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10635__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_255_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14709_ game.CPU.randy.counter1.count1\[2\] game.CPU.randy.counter1.count1\[1\] vssd1
+ vssd1 vccd1 vccd1 _08547_ sky130_fd_sc_hd__nand2_1
XANTENNA__09679__B game.CPU.applesa.ab.absxs.body_x\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15689_ _03225_ net352 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__xnor2_1
X_18477_ net636 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_188_Left_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17428_ net1274 _02856_ _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__a21o_1
XANTENNA__16771__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_177_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10618__B _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13585__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19699__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17359_ _02788_ net1114 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__and2b_1
XANTENNA__18073__A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13929__B game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_302_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16305__B _02303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload40 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__inv_8
XANTENNA_clkload48_A clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload51 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload51/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_301_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19029_ net1195 _00259_ _00700_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[74\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkload62 clknet_leaf_49_clk vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__inv_12
XANTENNA__14106__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout109_A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17079__A1 _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17079__B2 game.writer.tracker.frame\[393\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_266_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11449__B net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16826__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14117__A2_N net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11363__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_197_Left_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08994_ game.CPU.applesa.ab.absxs.body_x\[39\] vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__inv_2
XANTENNA__15663__A1_N net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1018_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19079__CLK net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout380_A _06209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16040__B net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_317_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11465__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09615_ net1086 game.CPU.applesa.ab.check_walls.above.walls\[3\] vssd1 vssd1 vccd1
+ vccd1 _03858_ sky130_fd_sc_hd__xor2_1
XANTENNA__11184__B net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16054__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12995__S net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_355_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13499__S0 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout645_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18248__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ net1102 game.CPU.applesa.ab.absxs.body_x\[113\] vssd1 vssd1 vccd1 vccd1 _03789_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_203_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17003__A1 _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_277_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14495__B _08368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09477_ net1156 net784 vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__or2_1
XANTENNA__18916__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09492__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16357__A3 _02341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16211__C1 _01838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09492__B2 net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16762__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload1 clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__inv_6
XFILLER_0_135_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16055__X _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ game.CPU.applesa.ab.check_walls.above.walls\[32\] net778 vssd1 vssd1 vccd1
+ vccd1 _05259_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_278_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16215__B net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13328__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_332_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10321_ net1439 _04501_ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_308_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14016__A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13423__S0 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13879__B2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_265_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13040_ net679 _06886_ _06913_ net504 vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__o211a_1
XFILLER_0_237_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10252_ _03493_ net747 vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_150_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10183_ net1125 _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout81_X net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1203 net1205 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16231__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1214 net1215 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08949__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1225 net1227 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__clkbuf_2
Xfanout1236 net1257 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__buf_2
X_14991_ net1227 net1254 game.CPU.applesa.ab.check_walls.above.walls\[19\] vssd1 vssd1
+ vccd1 vccd1 _00207_ sky130_fd_sc_hd__and3_1
Xfanout1247 net1257 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1258 game.CPU.kyle.L1.nextState\[1\] vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__clkbuf_4
Xfanout260 net262 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_4
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_4
Xfanout1269 game.CPU.applesa.ab.absxs.body_x\[49\] vssd1 vssd1 vccd1 vccd1 net1269
+ sky130_fd_sc_hd__buf_2
Xfanout282 net287 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_4
XFILLER_0_227_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16730_ net244 net172 _02320_ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__or3_2
X_13942_ net1075 game.CPU.applesa.ab.check_walls.above.walls\[64\] vssd1 vssd1 vccd1
+ vccd1 _07816_ sky130_fd_sc_hd__xor2_1
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__buf_2
XANTENNA__10314__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16045__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16661_ net153 net127 _02424_ _02548_ game.writer.tracker.frame\[123\] vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.next_frame\[123\] sky130_fd_sc_hd__a32o_1
XANTENNA__11094__B net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13873_ net1045 game.CPU.applesa.ab.check_walls.above.walls\[107\] vssd1 vssd1 vccd1
+ vccd1 _07747_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15253__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_319_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18400_ net617 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__inv_2
X_15612_ game.CPU.applesa.ab.absxs.body_x\[35\] net458 vssd1 vssd1 vccd1 vccd1 _01624_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12824_ game.writer.tracker.frame\[354\] game.writer.tracker.frame\[355\] net1001
+ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16592_ _02392_ _02493_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__nor2_1
X_19380_ clknet_leaf_3_clk _01386_ _00960_ vssd1 vssd1 vccd1 vccd1 game.CPU.bodymain1.main.score\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_15543_ net1066 _06551_ _01555_ _01563_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__a211o_1
XANTENNA__10617__A1 game.CPU.applesa.ab.absxs.body_x\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18331_ net616 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__inv_2
XANTENNA__18596__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12755_ game.writer.tracker.frame\[106\] game.writer.tracker.frame\[107\] net989
+ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__mux2_1
XANTENNA__09499__B net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19050__Q game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09483__A1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19841__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16821__A2_N net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09483__B2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11706_ game.CPU.applesa.ab.check_walls.above.walls\[165\] net315 _05592_ _05594_
+ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__a211o_1
X_18262_ net650 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__inv_2
X_15474_ _01470_ _01480_ _01492_ _01500_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_126_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16753__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12686_ net1076 net954 vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__nand2_4
XFILLER_0_194_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17213_ _02377_ net142 net119 _02734_ game.writer.tracker.frame\[489\] vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.next_frame\[489\] sky130_fd_sc_hd__a32o_1
X_14425_ _08297_ _08298_ vssd1 vssd1 vccd1 vccd1 _08299_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11637_ game.CPU.applesa.ab.check_walls.above.walls\[153\] net769 vssd1 vssd1 vccd1
+ vccd1 _05526_ sky130_fd_sc_hd__xor2_1
X_18193_ net612 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_210_Left_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17144_ net169 net69 net60 _02715_ net1636 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[439\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_315_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14356_ _08227_ _08228_ _08229_ vssd1 vssd1 vccd1 vccd1 _08230_ sky130_fd_sc_hd__and3_1
XANTENNA__16505__B1 _02449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_250_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11568_ game.CPU.applesa.ab.check_walls.above.walls\[128\] net773 vssd1 vssd1 vccd1
+ vccd1 _05457_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19991__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17702__C1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13307_ net505 _07178_ _07180_ net205 vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17075_ _02460_ net59 _02695_ net1713 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[390\]
+ sky130_fd_sc_hd__a22o_1
X_10519_ game.CPU.applesa.ab.absxs.body_x\[63\] net425 _04633_ net934 vssd1 vssd1
+ vccd1 vccd1 _01182_ sky130_fd_sc_hd__a22o_1
X_14287_ _03234_ net1069 net856 game.CPU.applesa.ab.absxs.body_y\[87\] vssd1 vssd1
+ vccd1 vccd1 _08161_ sky130_fd_sc_hd__o22a_1
XANTENNA__10454__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11499_ game.CPU.applesa.ab.check_walls.above.walls\[171\] net761 vssd1 vssd1 vccd1
+ vccd1 _05388_ sky130_fd_sc_hd__xor2_2
XANTENNA__16520__A3 _02460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_343_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire181_A _06638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16026_ _03228_ net343 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__xnor2_1
X_13238_ game.writer.tracker.frame\[478\] game.writer.tracker.frame\[479\] net1013
+ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__mux2_1
XANTENNA__19221__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11345__A2 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16808__A1 _02494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13169_ net512 _07042_ _07041_ net214 vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16141__A game.CPU.applesa.ab.absxs.body_x\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_236_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17977_ net590 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__inv_2
X_19716_ clknet_leaf_35_clk game.writer.tracker.next_frame\[311\] net1340 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[311\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_224_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15980__A game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16928_ net56 _02643_ _02650_ game.writer.tracker.frame\[288\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[288\] sky130_fd_sc_hd__a22o_1
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_284_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19371__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17233__A1 _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19647_ clknet_leaf_20_clk game.writer.tracker.next_frame\[242\] net1317 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[242\] sky130_fd_sc_hd__dfrtp_1
X_16859_ net133 _02410_ net122 _02625_ net1493 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[244\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_179_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09400_ net916 game.CPU.applesa.ab.check_walls.above.walls\[89\] _03430_ net1139
+ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19578_ clknet_leaf_31_clk game.writer.tracker.next_frame\[173\] net1294 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[173\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15795__B2 game.CPU.applesa.ab.absxs.body_x\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_149_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09331_ net919 game.CPU.applesa.ab.absxs.body_x\[82\] _03328_ net1125 vssd1 vssd1
+ vccd1 vccd1 _03574_ sky130_fd_sc_hd__a22o_1
X_18529_ net587 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__inv_2
XANTENNA__10608__B2 game.CPU.applesa.ab.absxs.body_x\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09474__A1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09474__B2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09262_ game.CPU.randy.counter1.count1\[5\] vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__inv_2
XFILLER_0_334_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_303_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13558__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ net797 vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__inv_2
XANTENNA__13022__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout226_A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16316__A _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_278_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_214_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12563__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16035__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10364__A game.CPU.walls.rand_wall.input2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1135_A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_274_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout595_A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13730__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__X _05635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__B2 game.CPU.applesa.ab.absxs.body_y\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1302_A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16051__A game.CPU.applesa.ab.absxs.body_x\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19714__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_328_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold13 game.CPU.reset_button1.eD1.D vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 game.CPU.walls.abc.number\[4\] vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ game.CPU.applesa.ab.absxs.body_x\[4\] vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout762_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19135__Q game.CPU.applesa.ab.check_walls.above.walls\[180\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 game.CPU.applesa.normal1.number\[6\] vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 game.CPU.applesa.twomode.number\[5\] vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_282_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11195__A game.CPU.applesa.ab.absxs.body_y\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold57 game.CPU.applesa.ab.x_final\[2\] vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_279_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold68 game.CPU.applesa.ab.absxs.body_y\[3\] vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 game.writer.tracker.frame\[237\] vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17224__A1 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout550_X net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1292_X net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19864__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10870_ _04751_ _04753_ _04763_ _04772_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__nand4_1
XFILLER_0_329_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13797__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11642__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09529_ net1089 _03445_ _03446_ net1135 _03769_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ game.CPU.applesa.ab.absxs.body_x\[41\] net377 net526 game.CPU.applesa.ab.absxs.body_y\[41\]
+ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_213_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10258__B net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_314_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12471_ _06347_ _06341_ _06346_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__or3b_1
XFILLER_0_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16226__A net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_352_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14210_ game.CPU.applesa.ab.absxs.body_x\[92\] net1070 vssd1 vssd1 vccd1 vccd1 _08084_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_193_Right_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15130__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11422_ _05300_ _05308_ _05309_ _05310_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__or4_1
X_15190_ _00018_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__inv_2
XFILLER_0_312_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12473__B net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14141_ _07842_ _07953_ _07973_ _08014_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__nand4_2
XFILLER_0_104_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_340_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11353_ game.CPU.applesa.ab.check_walls.above.walls\[136\] net773 vssd1 vssd1 vccd1
+ vccd1 _05242_ sky130_fd_sc_hd__xor2_1
XANTENNA__17160__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10304_ _04338_ net740 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__and2_2
XANTENNA__11089__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14072_ _07944_ _07945_ _07941_ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_293_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_265_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11284_ _04936_ _04938_ _05164_ _05173_ _05057_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__o311a_1
XANTENNA__15784__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11327__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13721__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13023_ _06864_ _06883_ net697 vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__mux2_1
X_17900_ net639 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__inv_2
X_10235_ _04424_ _04427_ _04426_ _04419_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09782__B game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18880_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[10\] _00575_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[10\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10535__B1 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1000 net1009 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__buf_2
Xfanout1011 net1013 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_280_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1022 net1041 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__buf_2
X_17831_ game.writer.updater.commands.count\[5\] _03158_ vssd1 vssd1 vccd1 vccd1 _03161_
+ sky130_fd_sc_hd__and2_1
Xfanout1033 net1034 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_280_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10166_ _04357_ _04360_ _04342_ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__o21a_1
XFILLER_0_218_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1044 net1051 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_8
Xfanout1055 net1059 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_163_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1066 net1068 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__buf_2
Xfanout1077 game.CPU.applesa.x\[0\] vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_4
X_17762_ _03109_ _03115_ _03117_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__and3_1
X_14974_ net1225 net1252 game.CPU.applesa.ab.check_walls.above.walls\[2\] vssd1 vssd1
+ vccd1 vccd1 _00099_ sky130_fd_sc_hd__and3_1
X_10097_ game.CPU.luck1.Qa\[0\] _04304_ net1162 vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__or3b_1
XANTENNA__15008__C net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1088 game.CPU.applesa.ab.snake_head_x\[3\] vssd1 vssd1 vccd1 vccd1 net1088
+ sky130_fd_sc_hd__buf_6
X_19501_ clknet_leaf_26_clk game.writer.tracker.next_frame\[96\] net1312 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[96\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17215__A1 _02299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1099 game.CPU.applesa.ab.snake_head_x\[1\] vssd1 vssd1 vccd1 vccd1 net1099
+ sky130_fd_sc_hd__buf_4
X_16713_ _02497_ net63 _02570_ net1655 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[152\]
+ sky130_fd_sc_hd__a22o_1
X_13925_ _07796_ _07797_ _07798_ _07788_ vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__o31a_1
XANTENNA__14029__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17693_ game.CPU.walls.rand_wall.count_luck\[7\] game.CPU.walls.rand_wall.count_luck\[6\]
+ _03071_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__and3_1
XANTENNA__14029__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload4_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19432_ clknet_leaf_39_clk game.writer.tracker.next_frame\[27\] net1352 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[27\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11833__A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16644_ net149 _02404_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__and2_1
X_13856_ net506 _07727_ _07728_ _07729_ net248 vssd1 vssd1 vccd1 vccd1 _07730_ sky130_fd_sc_hd__o221a_1
XFILLER_0_347_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13788__A0 game.writer.tracker.frame\[393\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12807_ game.writer.tracker.frame\[334\] game.writer.tracker.frame\[335\] net999
+ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__mux2_1
XANTENNA__09303__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__B net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19363_ clknet_leaf_69_clk _01369_ _00944_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16575_ net150 net127 _02497_ _02495_ net1543 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[88\]
+ sky130_fd_sc_hd__a32o_1
X_13787_ game.writer.tracker.frame\[397\] game.writer.tracker.frame\[399\] game.writer.tracker.frame\[400\]
+ game.writer.tracker.frame\[398\] net977 net1022 vssd1 vssd1 vccd1 vccd1 _07661_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09456__B2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10999_ game.CPU.applesa.ab.absxs.body_y\[47\] net399 vssd1 vssd1 vccd1 vccd1 _04889_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_270_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_252_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18314_ net620 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__inv_2
X_12738_ game.writer.tracker.frame\[68\] game.writer.tracker.frame\[69\] net1026 vssd1
+ vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__mux2_1
X_15526_ net1076 net1065 net1058 net1048 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16726__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15959__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19294_ clknet_leaf_69_clk _01338_ _00913_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.start_enable
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11263__B2 game.CPU.applesa.ab.absxs.body_y\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_270_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16407__Y _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15457_ _01450_ _01454_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__nand2_1
X_18245_ net644 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
XFILLER_0_316_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12669_ game.writer.updater.commands.mode\[1\] game.writer.updater.commands.mode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11015__A1 game.CPU.applesa.ab.absxs.body_x\[54\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14408_ game.CPU.applesa.ab.absxs.body_x\[44\] net890 net873 game.CPU.applesa.ab.absxs.body_x\[47\]
+ vssd1 vssd1 vccd1 vccd1 _08282_ sky130_fd_sc_hd__o22a_1
XANTENNA__11015__B2 game.CPU.applesa.ab.absxs.body_x\[55\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15388_ _08929_ vssd1 vssd1 vccd1 vccd1 _08930_ sky130_fd_sc_hd__inv_2
X_18176_ net608 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12383__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17127_ _02299_ net165 net76 _02710_ net1594 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[427\]
+ sky130_fd_sc_hd__a32o_1
X_14339_ _08211_ _08212_ vssd1 vssd1 vccd1 vccd1 _08213_ sky130_fd_sc_hd__nand2_1
Xhold505 game.writer.tracker.frame\[536\] vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10184__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold516 game.writer.tracker.frame\[126\] vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18351__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold527 game.CPU.applesa.ab.count_luck\[7\] vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 game.writer.tracker.frame\[103\] vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
X_17058_ _02592_ _02670_ net729 vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__o21a_1
XANTENNA__19737__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09973__A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold549 game.writer.tracker.frame\[155\] vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_284_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14504__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15694__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16009_ _03305_ net334 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19627__RESET_B net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_263_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _03651_ _03652_ _03656_ _04097_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__o31a_1
XFILLER_0_295_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14268__A1 game.CPU.applesa.ab.absxs.body_x\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18761__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14103__B net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19887__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13942__B game.CPU.applesa.ab.check_walls.above.walls\[64\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09695__A1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13434__S net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout176_A _06700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09695__B2 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11743__A game.CPU.applesa.ab.check_walls.above.walls\[157\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13228__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_295_Right_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_352_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_200_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11462__B net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09447__A1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_274_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09447__B2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_A game.CPU.walls.rand_wall.abduyd.next_wall\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1085_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09314_ net1094 game.CPU.applesa.ab.absxs.body_x\[66\] vssd1 vssd1 vccd1 vccd1 _03557_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_216_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17430__A net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15869__B net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19267__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09245_ net765 vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout510_A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_X net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13626__S0 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_X net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_322_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09176_ game.CPU.applesa.ab.check_walls.above.walls\[85\] vssd1 vssd1 vccd1 vccd1
+ _03425_ sky130_fd_sc_hd__inv_2
XFILLER_0_334_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12293__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_322_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17142__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18261__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1138_X net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18969__Q game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xoutput14 net14 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout977_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput36 net36 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_285_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_247_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10517__B1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_227_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout89_A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ net1081 _04224_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__or2_1
XANTENNA__11637__B net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13467__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout932_X net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ game.CPU.applesa.ab.apple_possible\[7\] _05193_ vssd1 vssd1 vccd1 vccd1 _05858_
+ sky130_fd_sc_hd__xor2_2
XFILLER_0_203_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_199_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20031__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09686__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13710_ game.writer.tracker.frame\[233\] game.writer.tracker.frame\[235\] game.writer.tracker.frame\[236\]
+ game.writer.tracker.frame\[234\] net968 net998 vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__mux4_1
XANTENNA__11653__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ net543 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.next_head\[5\] sky130_fd_sc_hd__clkinv_4
X_14690_ game.CPU.randy.counter1.count1\[15\] _08499_ _08500_ game.CPU.randy.counter1.count1\[13\]
+ _08528_ vssd1 vssd1 vccd1 vccd1 _08529_ sky130_fd_sc_hd__a221o_1
XANTENNA__16956__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_262_Right_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_316_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12468__B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13641_ game.writer.tracker.frame\[57\] game.writer.tracker.frame\[59\] game.writer.tracker.frame\[60\]
+ game.writer.tracker.frame\[58\] net980 net1040 vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_296_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09438__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10853_ game.CPU.randy.counter1.count1\[12\] _03501_ game.CPU.randy.counter1.count\[11\]
+ _03502_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_66_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09438__B2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_238_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16360_ net177 _02240_ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__nor2_1
X_13572_ game.writer.tracker.frame\[353\] game.writer.tracker.frame\[355\] game.writer.tracker.frame\[356\]
+ game.writer.tracker.frame\[354\] net976 net1009 vssd1 vssd1 vccd1 vccd1 _07446_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12442__B1 game.CPU.applesa.twoapples.absxs.next_head\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__B2 game.CPU.applesa.ab.absxs.body_y\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10784_ game.CPU.applesa.ab.absxs.body_y\[56\] net328 _04723_ net935 vssd1 vssd1
+ vccd1 vccd1 _01007_ sky130_fd_sc_hd__a22o_1
X_15311_ net757 _08854_ _08855_ _08856_ _08857_ vssd1 vssd1 vccd1 vccd1 _08858_ sky130_fd_sc_hd__a32o_1
XFILLER_0_183_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12523_ game.CPU.applesa.ab.absxs.body_x\[71\] net530 vssd1 vssd1 vccd1 vccd1 _06400_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16291_ net2041 net720 _02292_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[9\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__16184__A1 _02133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_313_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16723__A3 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15242_ net2036 _08802_ vssd1 vssd1 vccd1 vccd1 _08803_ sky130_fd_sc_hd__nand2_1
X_18030_ net590 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__inv_2
XANTENNA__14195__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12454_ game.CPU.applesa.ab.absxs.body_x\[51\] net531 net360 game.CPU.applesa.ab.absxs.body_y\[48\]
+ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11405_ net806 net316 net260 game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1
+ vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__o2bb2a_1
X_15173_ game.CPU.bodymain1.main.score\[7\] net1114 net1115 vssd1 vssd1 vccd1 vccd1
+ _08749_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12385_ game.CPU.applesa.ab.absxs.body_x\[27\] net529 vssd1 vssd1 vccd1 vccd1 _06262_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10756__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_327_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14124_ net956 game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1 vccd1
+ vccd1 _07998_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09793__A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11336_ game.CPU.applesa.ab.check_walls.above.walls\[80\] net775 vssd1 vssd1 vccd1
+ vccd1 _05225_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19981_ clknet_leaf_47_clk _01405_ net1298 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.y\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18784__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13519__S net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_249_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14055_ net983 net790 vssd1 vssd1 vccd1 vccd1 _07929_ sky130_fd_sc_hd__or2_1
X_18932_ clknet_leaf_5_clk net7 _00616_ vssd1 vssd1 vccd1 vccd1 game.CPU.start_pause_button1.sync1.Q
+ sky130_fd_sc_hd__dfrtp_1
X_11267_ _04856_ _04857_ _04859_ _04860_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a22o_1
XANTENNA__10508__B1 _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13170__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ game.writer.tracker.frame\[548\] game.writer.tracker.frame\[549\] net1006
+ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__mux2_1
X_10218_ _04409_ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__xnor2_1
X_18863_ clknet_leaf_1_clk _01254_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15019__B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11198_ _03316_ net404 vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__xnor2_1
X_17814_ game.writer.updater.commands.count\[0\] _03148_ vssd1 vssd1 vccd1 vccd1 _03149_
+ sky130_fd_sc_hd__nor2_1
X_10149_ game.CPU.randy.f1.state\[1\] game.CPU.randy.f1.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _04344_ sky130_fd_sc_hd__nand2b_2
X_18794_ clknet_leaf_9_clk _01209_ _00531_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17745_ _03360_ _03102_ _03106_ vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__a21oi_1
X_14957_ _08678_ _08681_ _08679_ _08661_ vssd1 vssd1 vccd1 vccd1 _08734_ sky130_fd_sc_hd__o211a_1
XANTENNA__19503__Q game.writer.tracker.frame\[98\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13107__X _06981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15035__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_338_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13908_ net938 game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1 vccd1
+ vccd1 _07782_ sky130_fd_sc_hd__xor2_1
X_17676_ _03523_ _03060_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__and2_1
X_14888_ _08663_ _08664_ vssd1 vssd1 vccd1 vccd1 _08665_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19415_ clknet_leaf_48_clk game.writer.tracker.next_frame\[10\] net1297 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[10\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16411__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09033__A game.CPU.applesa.ab.absxs.body_x\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16627_ _02377_ _02518_ _02532_ net1643 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[105\]
+ sky130_fd_sc_hd__a22o_1
X_13839_ _07711_ _07712_ net506 vssd1 vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__mux2_1
XANTENNA__09429__A1 game.CPU.applesa.ab.snake_head_x\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_328_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19346_ clknet_leaf_72_clk _01361_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.enablea2
+ sky130_fd_sc_hd__dfxtp_1
X_16558_ net222 _02407_ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__nor2_4
XANTENNA__15689__B net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12433__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15509_ net879 _06555_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19277_ clknet_leaf_7_clk _00047_ _00907_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_16489_ net168 net56 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__and2_2
XFILLER_0_72_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09030_ game.CPU.applesa.ab.absxs.body_x\[26\] vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__inv_2
XANTENNA__14186__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18228_ net665 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18159_ net635 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_349_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold302 game.CPU.randy.counter1.count\[13\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_211_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold313 game.writer.tracker.frame\[485\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 game.writer.tracker.frame\[58\] vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold335 game.CPU.randy.f1.a1.count\[3\] vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 game.writer.tracker.frame\[514\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload30_A clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold357 game.writer.tracker.frame\[317\] vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_257_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10913__Y game.CPU.applesa.ab.absxs.next_head\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold368 game.CPU.kyle.L1.cnt_500hz\[11\] vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09932_ _04158_ _04169_ _04170_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__and3_1
Xhold379 game.writer.tracker.frame\[106\] vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout804 game.CPU.applesa.ab.check_walls.above.walls\[101\] vssd1 vssd1 vccd1 vccd1
+ net804 sky130_fd_sc_hd__buf_2
XFILLER_0_256_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout815 game.CPU.applesa.ab.check_walls.above.walls\[69\] vssd1 vssd1 vccd1 vccd1
+ net815 sky130_fd_sc_hd__clkbuf_4
X_20052_ net1370 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
Xfanout826 game.CPU.applesa.ab.check_walls.above.walls\[28\] vssd1 vssd1 vccd1 vccd1
+ net826 sky130_fd_sc_hd__clkbuf_4
Xfanout837 net839 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_4
XFILLER_0_272_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09863_ net905 game.CPU.applesa.ab.absxs.body_y\[46\] _03310_ net1150 vssd1 vssd1
+ vccd1 vccd1 _04106_ sky130_fd_sc_hd__a22o_1
Xfanout848 net849 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__clkbuf_4
Xfanout859 net860 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_175_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13449__C1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1000_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09794_ net926 game.CPU.applesa.ab.absxs.body_x\[43\] game.CPU.applesa.ab.absxs.body_x\[41\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_300_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16650__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout460_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_222_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11473__A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14487__C _08359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12288__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout725_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_327_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13847__S0 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18256__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14413__B2 game.CPU.applesa.ab.absxs.body_y\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_X net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18657__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19902__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09597__B game.CPU.applesa.ab.absxs.body_x\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09840__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1255_X net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16705__A3 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09840__B2 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_311_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14177__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09228_ game.CPU.applesa.ab.check_walls.above.walls\[179\] vssd1 vssd1 vccd1 vccd1
+ _03477_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_233_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09159_ game.CPU.applesa.ab.check_walls.above.walls\[51\] vssd1 vssd1 vccd1 vccd1
+ _03408_ sky130_fd_sc_hd__inv_2
XFILLER_0_310_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12170_ net788 net293 net288 game.CPU.applesa.ab.check_walls.above.walls\[158\] vssd1
+ vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__18699__Q game.CPU.applesa.ab.absxs.body_x\[49\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_248_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17130__A3 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13339__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11950__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ _03353_ net404 vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_287_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13152__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_331_Right_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11052_ _03321_ net536 vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10271__B game.CPU.applesa.ab.apple_possible\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11163__B1 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10003_ net914 _04210_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_322_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ game.CPU.applesa.ab.absxs.body_y\[115\] net435 vssd1 vssd1 vccd1 vccd1 _01872_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_262_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14811_ game.CPU.randy.counter1.count\[12\] _08619_ vssd1 vssd1 vccd1 vccd1 _08621_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_188_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12479__A game.CPU.applesa.ab.absxs.body_x\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15791_ _01794_ _01795_ _01799_ _01800_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__or4_1
XANTENNA__13455__A2 _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19432__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17530_ game.CPU.kyle.L1.row_2\[72\] _02774_ net428 vssd1 vssd1 vccd1 vccd1 _02958_
+ sky130_fd_sc_hd__and3_1
X_11954_ game.CPU.applesa.ab.check_walls.above.walls\[118\] net299 _05840_ _05841_
+ _05833_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__o221a_1
XFILLER_0_98_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14742_ game.CPU.randy.counter1.count1\[13\] _08567_ vssd1 vssd1 vccd1 vccd1 _08569_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__16929__B1 _02650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12198__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10905_ game.CPU.applesa.ab.check_walls.collision_left _04802_ _04803_ _04806_ vssd1
+ vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_86_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17461_ _02888_ _02889_ _02785_ _02789_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__o211ai_2
X_14673_ game.CPU.randy.counter1.count1\[4\] _04347_ _08501_ game.CPU.randy.counter1.count1\[5\]
+ vssd1 vssd1 vccd1 vccd1 _08512_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ net827 net312 vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__nand2_1
XFILLER_0_168_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13838__S0 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_317_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19200_ clknet_leaf_67_clk _01309_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13624_ _07496_ _07497_ net512 vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__mux2_1
X_16412_ net196 _02340_ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__or2_2
XFILLER_0_345_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10836_ game.CPU.randy.counter1.count\[17\] _03496_ game.CPU.randy.counter1.count\[16\]
+ _03497_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__o22a_1
XANTENNA__19582__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17392_ _02783_ _02820_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__or2_1
XFILLER_0_345_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19131_ net1184 _00172_ _00802_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[176\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12966__B2 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13555_ _07427_ _07428_ net488 vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__mux2_2
X_16343_ net197 _02330_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__nor2_2
XFILLER_0_27_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_333_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10767_ game.CPU.applesa.ab.absxs.body_y\[81\] _04673_ _04674_ game.CPU.applesa.ab.absxs.body_y\[77\]
+ vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__a22o_1
X_12506_ _03332_ net369 vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_171_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16274_ _02245_ net236 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__nor2_2
X_19062_ net1191 _00096_ _00733_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[107\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10441__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ net502 _07136_ _07359_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15021__C game.CPU.applesa.ab.check_walls.above.walls\[49\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ game.CPU.applesa.ab.absxs.body_y\[84\] _04610_ _04611_ game.CPU.applesa.ab.absxs.body_y\[80\]
+ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10446__B net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15225_ game.CPU.applesa.normal1.number\[1\] _08785_ vssd1 vssd1 vccd1 vccd1 _08790_
+ sky130_fd_sc_hd__or2_1
X_18013_ net639 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__inv_2
XFILLER_0_340_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12437_ game.CPU.applesa.ab.absxs.body_y\[105\] net524 vssd1 vssd1 vccd1 vccd1 _06314_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_313_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16414__A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_340_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15156_ net1213 net1240 game.CPU.applesa.ab.check_walls.above.walls\[184\] vssd1
+ vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__and3_1
X_12368_ game.CPU.applesa.ab.absxs.body_y\[6\] net519 vssd1 vssd1 vccd1 vccd1 _06245_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_266_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14107_ net878 game.CPU.applesa.ab.check_walls.above.walls\[50\] game.CPU.applesa.ab.check_walls.above.walls\[51\]
+ net875 _07976_ vssd1 vssd1 vccd1 vccd1 _07981_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_39_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11319_ net814 net256 _05205_ _05203_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__o211a_1
X_19964_ clknet_leaf_44_clk game.writer.tracker.next_frame\[559\] net1306 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[559\] sky130_fd_sc_hd__dfrtp_1
X_15087_ net1206 net1243 game.CPU.applesa.ab.check_walls.above.walls\[115\] vssd1
+ vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__and3_1
XFILLER_0_293_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12299_ net827 _04782_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_52_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_160_Left_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14038_ net983 net799 vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__xnor2_1
X_18915_ clknet_leaf_4_clk net1401 _00599_ vssd1 vssd1 vccd1 vccd1 game.CPU.up_button.eD1.Q2
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15972__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19895_ clknet_leaf_14_clk game.writer.tracker.next_frame\[490\] net1287 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[490\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09898__A1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18846_ clknet_leaf_0_clk _01237_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16632__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_350_Left_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18777_ clknet_leaf_64_clk _01194_ _00514_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[87\]
+ sky130_fd_sc_hd__dfrtp_4
X_15989_ _01997_ _01998_ _01999_ _02000_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a22o_1
X_17728_ net2015 _03093_ _03095_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_292_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19925__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17659_ game.CPU.kyle.L1.cnt_500hz\[9\] game.CPU.kyle.L1.cnt_500hz\[10\] _03047_
+ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__and3_1
XFILLER_0_309_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_258_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18076__A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_271_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16308__B net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19329_ clknet_leaf_72_clk net1417 _00934_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twomode.number\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_193_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14159__B1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_311_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ game.CPU.applesa.ab.absxs.body_x\[96\] vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__inv_2
XANTENNA__13948__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout306_A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13382__A1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1048_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19305__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_304_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold110 game.writer.tracker.frame\[494\] vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 game.writer.tracker.frame\[350\] vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 game.writer.tracker.frame\[482\] vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 game.writer.tracker.frame\[402\] vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16043__B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold154 game.writer.tracker.frame\[574\] vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_269_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold165 game.writer.tracker.frame\[268\] vssd1 vssd1 vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 game.CPU.randy.f1.c1.count\[13\] vssd1 vssd1 vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_282_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1215_A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 game.writer.tracker.frame\[43\] vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 net604 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__buf_4
Xhold198 game.writer.tracker.frame\[238\] vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 net624 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14331__B1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16871__A2 _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11187__B net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15882__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09915_ game.CPU.applesa.clk_body game.CPU.bodymain1.main.pause_clk vssd1 vssd1 vccd1
+ vccd1 _04157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_229_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout623 net624 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__buf_2
Xfanout634 net651 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_4
XANTENNA_fanout675_A _07401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19455__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_298_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout296_X net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 net646 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_4
Xfanout656 net657 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__buf_4
XFILLER_0_186_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout667 net670 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_2
X_20035_ net1383 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
X_09846_ net1090 game.CPU.applesa.ab.absxs.body_x\[30\] vssd1 vssd1 vccd1 vccd1 _04089_
+ sky130_fd_sc_hd__xor2_1
Xfanout678 net681 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_4
Xfanout689 net691 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_336_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09777_ net1082 game.CPU.applesa.ab.check_walls.above.walls\[147\] vssd1 vssd1 vccd1
+ vccd1 _04020_ sky130_fd_sc_hd__xor2_1
XANTENNA__13437__A2 _06956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout842_A _06574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12299__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16994__A _02455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12645__B1 _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09340__A2_N net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18982__Q game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10120__A1 game.CPU.applesa.enable_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16058__X _02070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_293_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ net794 net254 net249 game.CPU.applesa.ab.check_walls.above.walls\[124\] _05558_
+ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__a221o_1
XFILLER_0_352_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_235_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12948__A1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16218__B net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10621_ net1080 _04679_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__nor2_2
XANTENNA__09813__A1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09813__B2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13340_ net219 _07213_ net276 vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__a21o_1
XANTENNA__09895__X _04138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10552_ game.CPU.applesa.ab.absxs.body_x\[30\] net330 _04649_ net930 vssd1 vssd1
+ vccd1 vccd1 _01165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_322_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ game.writer.tracker.frame\[492\] game.writer.tracker.frame\[493\] net995
+ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__mux2_1
X_10483_ _04583_ _04591_ _04606_ net850 vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__a211o_4
XANTENNA__16234__A _02237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_297_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15010_ net1215 net1241 net822 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__and3_1
XANTENNA__13373__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12222_ net811 net423 vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_350_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17103__A3 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11378__A game.CPU.applesa.ab.check_walls.above.walls\[179\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_248_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ game.CPU.applesa.ab.check_walls.above.walls\[135\] net293 vssd1 vssd1 vccd1
+ vccd1 _06040_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09119__Y _03368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16521__X _02461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16888__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_246_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11104_ game.CPU.applesa.ab.absxs.body_x\[35\] net408 vssd1 vssd1 vccd1 vccd1 _04994_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__11097__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16961_ _02418_ net94 _02659_ net1857 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[312\]
+ sky130_fd_sc_hd__a22o_1
X_12084_ game.CPU.applesa.ab.check_walls.above.walls\[20\] net554 vssd1 vssd1 vccd1
+ vccd1 _05971_ sky130_fd_sc_hd__or2_1
XANTENNA__13676__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18700_ clknet_leaf_12_clk _01117_ _00437_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[50\]
+ sky130_fd_sc_hd__dfrtp_4
X_11035_ game.CPU.applesa.ab.absxs.body_x\[65\] net412 net401 _03334_ vssd1 vssd1
+ vccd1 vccd1 _04925_ sky130_fd_sc_hd__a22o_1
X_15912_ _03447_ net354 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__nand2_1
X_19680_ clknet_leaf_34_clk game.writer.tracker.next_frame\[275\] net1322 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[275\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11687__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16892_ net200 net68 net93 _02639_ net1483 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[263\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__11687__B2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19948__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18631_ clknet_leaf_10_clk _01048_ _00368_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11825__B net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15843_ net828 net442 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19053__Q game.CPU.applesa.ab.check_walls.above.walls\[98\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15822__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18562_ clknet_leaf_9_clk _00982_ _00299_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_12986_ net183 net174 vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__nand2_1
X_15774_ _01782_ _01783_ _01784_ _01785_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__or4_1
XFILLER_0_204_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12002__A game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17513_ net1454 net264 _02880_ _02941_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_335_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14725_ game.CPU.randy.counter1.count1\[7\] _08555_ vssd1 vssd1 vccd1 vccd1 _08558_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_358_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11937_ net572 _05589_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ net617 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__inv_2
XANTENNA__14389__B1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17444_ _02825_ _02847_ _02873_ _03218_ _02773_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_262_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10662__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11868_ net574 _05399_ _05402_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__a21oi_1
X_14656_ game.CPU.randy.counter1.count1\[17\] _08492_ _08494_ game.CPU.randy.counter1.count1\[16\]
+ vssd1 vssd1 vccd1 vccd1 _08495_ sky130_fd_sc_hd__o22ai_1
XANTENNA__12939__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13607_ game.writer.tracker.frame\[293\] game.writer.tracker.frame\[295\] game.writer.tracker.frame\[296\]
+ game.writer.tracker.frame\[294\] net964 net988 vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__mux4_1
XANTENNA__11560__B _05213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ game.CPU.applesa.ab.absxs.body_y\[10\] _04689_ _04707_ game.CPU.applesa.ab.absxs.body_y\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17375_ net1117 _02802_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__nand2_1
X_14587_ net1275 _03521_ _08448_ game.CPU.clock1.counter\[15\] game.CPU.clock1.counter\[19\]
+ vssd1 vssd1 vccd1 vccd1 _08449_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11799_ game.CPU.applesa.ab.check_walls.above.walls\[196\] net392 net307 game.CPU.applesa.ab.check_walls.above.walls\[197\]
+ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_156_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_305_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19114_ net1181 _00153_ _00785_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[159\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__19328__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16326_ game.writer.tracker.frame\[17\] net722 _02312_ _02319_ net136 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.next_frame\[17\] sky130_fd_sc_hd__a32o_1
X_13538_ _07410_ _07411_ net493 vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__mux2_1
XANTENNA__15967__B net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10176__B game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_298_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19045_ net1192 _00277_ _00716_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[90\]
+ sky130_fd_sc_hd__dfrtp_4
X_13469_ net512 _07087_ _07342_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__o21ai_1
X_16257_ _02245_ _02262_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_301_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15208_ game.CPU.applesa.normal1.number\[6\] _08770_ game.CPU.applesa.normal1.counter
+ vssd1 vssd1 vccd1 vccd1 _08776_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_346_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_313_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10178__A1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16188_ _02158_ _02199_ _02159_ _02197_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__or4b_4
XANTENNA__12391__B net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19478__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10192__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15139_ net1210 net1236 net786 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__and3_1
XANTENNA__16431__X _02394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_266_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_294_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19947_ clknet_leaf_38_clk game.writer.tracker.next_frame\[542\] net1324 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[542\] sky130_fd_sc_hd__dfrtp_1
X_09700_ net904 game.CPU.applesa.ab.check_walls.above.walls\[62\] net816 net908 vssd1
+ vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__a22o_1
XFILLER_0_281_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19878_ clknet_leaf_27_clk game.writer.tracker.next_frame\[473\] net1316 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[473\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10920__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17802__A1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11405__A2_N net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ net1092 game.CPU.applesa.ab.absxs.body_x\[18\] vssd1 vssd1 vccd1 vccd1 _03874_
+ sky130_fd_sc_hd__xor2_1
X_18829_ clknet_leaf_3_clk _01220_ _00557_ vssd1 vssd1 vccd1 vccd1 game.CPU.bodymain1.Direction\[0\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__17802__B2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14111__B game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15813__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ net927 game.CPU.applesa.ab.absxs.body_x\[63\] game.CPU.applesa.ab.absxs.body_y\[63\]
+ net908 _03804_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__a221o_1
XANTENNA__12627__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13824__C1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10102__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09493_ _03728_ _03729_ _03731_ _03732_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__or4_1
XANTENNA__10102__B2 net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11751__A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17030__A2 _02670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10653__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11850__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16038__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout423_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11602__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout211_X net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16541__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12582__A game.CPU.applesa.ab.absxs.body_x\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1332_A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_230_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13355__B2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout792_A game.CPU.applesa.ab.check_walls.above.walls\[133\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__B _04702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15893__A game.CPU.applesa.ab.absxs.body_x\[40\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13107__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1218_X net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14304__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout420 _04784_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13658__A2 game.writer.tracker.frame\[48\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout431 net437 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13617__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout442 net443 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_4
XANTENNA__11669__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout453 net454 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout71_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout464 _08423_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_4
XANTENNA__14302__A game.CPU.applesa.ab.absxs.body_y\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16995__Y _02670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_272_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout475 _08418_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_4
XANTENNA__16057__B1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout486 _06596_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_2
X_20018_ net1276 vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xfanout497 net499 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_4
X_09829_ net908 game.CPU.applesa.ab.absxs.body_y\[15\] game.CPU.applesa.ab.absxs.body_y\[13\]
+ net899 _04065_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__a221o_1
XANTENNA__11645__B _05504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18995__CLK net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ game.writer.tracker.frame\[280\] game.writer.tracker.frame\[281\] net1018
+ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_241_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12618__B1 game.CPU.applesa.twoapples.absxs.next_head\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12771_ game.writer.tracker.frame\[84\] game.writer.tracker.frame\[85\] net1029 vssd1
+ vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__mux2_1
XANTENNA__10829__X _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16229__A net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13830__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17021__A2 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15133__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14510_ game.CPU.apple_location2\[0\] net886 net938 _03203_ vssd1 vssd1 vccd1 vccd1
+ _08384_ sky130_fd_sc_hd__a22o_1
X_11722_ game.CPU.applesa.ab.check_walls.above.walls\[76\] net395 _05609_ vssd1 vssd1
+ vccd1 vccd1 _05610_ sky130_fd_sc_hd__o21ba_1
X_15490_ _01513_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__inv_2
XANTENNA__11841__A1 game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12476__B net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__A game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19564__RESET_B net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14441_ game.CPU.applesa.ab.absxs.body_x\[90\] net1053 vssd1 vssd1 vccd1 vccd1 _08315_
+ sky130_fd_sc_hd__nand2_1
X_11653_ net567 _05540_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__nor2_1
XANTENNA__16780__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16516__X _02458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout60 _02692_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_4
XANTENNA__18444__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15583__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout71 net72 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_4
X_10604_ game.CPU.applesa.ab.absxs.body_x\[89\] _04590_ net329 game.CPU.applesa.ab.absxs.body_x\[85\]
+ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_155_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout82 _02690_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__buf_4
X_17160_ _02444_ _02719_ net558 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__a21oi_1
X_14372_ game.CPU.applesa.ab.absxs.body_x\[116\] net889 net985 _03355_ vssd1 vssd1
+ vccd1 vccd1 _08246_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_330_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout93 net97 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_2
XFILLER_0_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ _05391_ _05394_ _05408_ _05472_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15787__B net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16235__Y _02243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ net688 _06713_ _07196_ net229 vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__o211a_1
X_16111_ game.CPU.applesa.ab.absxs.body_x\[57\] net473 net441 game.CPU.applesa.ab.absxs.body_y\[58\]
+ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10535_ game.CPU.applesa.ab.absxs.body_x\[47\] _04640_ _04641_ game.CPU.applesa.ab.absxs.body_x\[43\]
+ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__a22o_1
X_17091_ _02484_ net58 _02699_ net1528 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[402\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19620__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13346__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13254_ net226 _07127_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__or2_1
X_16042_ game.CPU.applesa.ab.absxs.body_y\[44\] net341 vssd1 vssd1 vccd1 vccd1 _02054_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10466_ net931 game.CPU.applesa.ab.absxs.body_x\[97\] _04594_ _04598_ vssd1 vssd1
+ vccd1 vccd1 _01200_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19048__Q game.CPU.applesa.ab.check_walls.above.walls\[93\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12205_ _06083_ _06085_ _06086_ _06087_ _06090_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__o32a_1
XFILLER_0_122_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17088__A2 _02692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ net217 _07052_ _07058_ net285 vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__o211a_1
X_10397_ _03220_ game.CPU.randy.f1.state\[4\] _04547_ _04360_ vssd1 vssd1 vccd1 vccd1
+ _04548_ sky130_fd_sc_hd__a31o_1
X_19801_ clknet_leaf_33_clk game.writer.tracker.next_frame\[396\] net1324 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[396\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19770__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09970__B1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12136_ _05197_ _05199_ _05200_ _05202_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__or4_1
XANTENNA__17066__Y _02690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17993_ net656 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__inv_2
X_19732_ clknet_leaf_19_clk game.writer.tracker.next_frame\[327\] net1335 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[327\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11836__A game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16944_ game.writer.tracker.frame\[300\] _02654_ vssd1 vssd1 vccd1 vccd1 _02655_
+ sky130_fd_sc_hd__and2_1
X_12067_ net795 net386 vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_166_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10740__A game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_341_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output52_A net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09306__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ game.CPU.applesa.ab.absxs.body_x\[89\] net323 vssd1 vssd1 vccd1 vccd1 _04908_
+ sky130_fd_sc_hd__nand2_1
X_19663_ clknet_leaf_32_clk game.writer.tracker.next_frame\[258\] net1291 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[258\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11555__B net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16875_ _02552_ net107 _02630_ net1803 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[255\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19000__CLK net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18614_ clknet_leaf_13_clk _01031_ _00351_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[108\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17260__A2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15826_ _01828_ _01829_ _01835_ _01837_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__or4b_2
XANTENNA__12609__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19594_ clknet_leaf_36_clk game.writer.tracker.next_frame\[189\] net1355 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[189\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13806__C1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14074__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18545_ net632 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__inv_2
X_15757_ _03316_ net339 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__xnor2_1
X_12969_ net490 _06842_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__or2_1
XANTENNA__15043__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17012__A2 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14708_ game.CPU.randy.counter1.count1\[2\] game.CPU.randy.counter1.count1\[1\] vssd1
+ vssd1 vccd1 vccd1 _08546_ sky130_fd_sc_hd__or2_1
XANTENNA__19150__CLK net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10635__A2 game.CPU.applesa.ab.absxs.body_x\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_255_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11832__A1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18476_ net638 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15688_ game.CPU.applesa.ab.absxs.body_y\[6\] net440 vssd1 vssd1 vccd1 vccd1 _01700_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12386__B net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09041__A game.CPU.applesa.ab.absxs.body_x\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15978__A game.CPU.applesa.ab.check_walls.above.walls\[68\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18718__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17427_ _02783_ _02828_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14639_ game.CPU.clock1.counter\[19\] _08480_ net267 vssd1 vssd1 vccd1 vccd1 _08482_
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_103_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16771__A1 _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16426__X _02391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_14_clk_X clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17358_ net1115 net1114 game.CPU.bodymain1.main.score\[7\] vssd1 vssd1 vccd1 vccd1
+ _02788_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_119_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16309_ net971 _02246_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__nand2_1
XFILLER_0_302_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17289_ game.writer.tracker.frame\[546\] _02753_ vssd1 vssd1 vccd1 vccd1 _02754_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10915__A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload30 clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 clkload30/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload41 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload41/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_301_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19028_ net1193 _00258_ _00699_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[73\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkload52 clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload63 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__clkinv_8
XANTENNA_clkbuf_leaf_29_clk_X clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14106__B game.CPU.applesa.ab.check_walls.above.walls\[48\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11899__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_266_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_208_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08993_ game.CPU.applesa.ab.absxs.body_x\[47\] vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13196__S0 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10650__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_305_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout373_A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18529__A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ _03854_ _03855_ _03856_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__or3_1
XANTENNA__13499__S1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ net1093 game.CPU.applesa.ab.absxs.body_x\[114\] vssd1 vssd1 vccd1 vccd1 _03788_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_203_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout540_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11989__A2_N net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16049__A game.CPU.applesa.ab.absxs.body_y\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_333_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout638_A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_277_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09476_ net1156 net784 vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_290_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_219_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_309_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16211__B1 _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16762__A1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19643__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10097__A game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1070_X net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout805_A game.CPU.applesa.ab.check_walls.above.walls\[94\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18264__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload2 clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__inv_6
XFILLER_0_135_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_352_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13328__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10320_ game.CPU.randy.f1.a1.count\[12\] game.CPU.randy.f1.a1.count\[11\] _04500_
+ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__and3_1
XANTENNA__19793__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_308_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13423__S1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13695__X _07569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10251_ net767 _04441_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16817__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ net1168 game.CPU.applesa.ab.apple_possible\[7\] vssd1 vssd1 vccd1 vccd1 _04375_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout962_X net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10831__Y _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10562__A1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1204 net1205 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_243_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1215 net1216 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__buf_2
XFILLER_0_273_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1226 net1227 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__buf_1
XANTENNA__11656__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1237 net1242 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__clkbuf_2
Xfanout250 net251 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_2
X_14990_ net1223 net1250 game.CPU.applesa.ab.check_walls.above.walls\[18\] vssd1 vssd1
+ vccd1 vccd1 _00206_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout74_X net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1248 net1249 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13500__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1259 game.CPU.kyle.L1.nextState\[0\] vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__clkbuf_4
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09126__A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout272 net273 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_4
Xfanout283 net284 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_245_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20000__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13941_ net1058 game.CPU.applesa.ab.check_walls.above.walls\[66\] vssd1 vssd1 vccd1
+ vccd1 _07815_ sky130_fd_sc_hd__xor2_1
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_198_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16660_ _02243_ net157 _02425_ net731 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__o31a_1
XANTENNA__17242__A2 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19173__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13872_ net940 net800 vssd1 vssd1 vccd1 vccd1 _07746_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_260_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08965__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15611_ _01619_ _01620_ _01621_ _01622_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_319_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12823_ game.writer.tracker.frame\[360\] game.writer.tracker.frame\[361\] net1001
+ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__mux2_1
X_16591_ net1619 _02505_ _02507_ net126 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[94\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_201_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13803__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11391__A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18330_ net616 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__inv_2
X_15542_ net1066 net1049 net1057 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10617__A2 _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__Y _03381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12754_ game.writer.tracker.frame\[108\] game.writer.tracker.frame\[109\] net995
+ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__mux2_1
XANTENNA__09483__A2 game.CPU.applesa.ab.check_walls.above.walls\[177\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16202__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11705_ game.CPU.applesa.ab.check_walls.above.walls\[164\] net250 _05593_ vssd1 vssd1
+ vccd1 vccd1 _05594_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_139_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18261_ net650 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
XFILLER_0_343_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16753__A1 _02535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12685_ net943 _06556_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__xnor2_4
X_15473_ _01463_ _01482_ _01487_ _01499_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__o211ai_1
XANTENNA__13810__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17212_ _02530_ _02720_ net714 vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__o21a_1
X_14424_ _03258_ net1059 net994 _03324_ _08291_ vssd1 vssd1 vccd1 vccd1 _08298_ sky130_fd_sc_hd__o221a_1
X_11636_ net746 _05524_ _05523_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__o21ai_1
X_18192_ net609 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17143_ net166 _02415_ net81 _02715_ net1465 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[438\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__16505__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11567_ net792 net314 vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__nor2_1
X_14355_ _08221_ _08222_ _08223_ _08225_ vssd1 vssd1 vccd1 vccd1 _08229_ sky130_fd_sc_hd__and4_1
XFILLER_0_107_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16505__B2 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13306_ net481 _07179_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__or2_1
X_10518_ _03270_ _04632_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__nor2_1
X_17074_ _02456_ _02693_ net736 vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__o21a_1
XFILLER_0_296_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14286_ game.CPU.applesa.ab.absxs.body_x\[87\] net876 net861 game.CPU.applesa.ab.absxs.body_y\[85\]
+ _08159_ vssd1 vssd1 vccd1 vccd1 _08160_ sky130_fd_sc_hd__o221a_1
X_11498_ net746 _05385_ _05383_ _05382_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13237_ game.writer.tracker.frame\[474\] game.writer.tracker.frame\[475\] net1017
+ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_268_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16025_ _03229_ net347 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_343_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10449_ net1117 net1119 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16808__A2 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_268_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12542__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13168_ _07031_ _07033_ net689 vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_283_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16141__B net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13178__S0 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11566__A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ net785 net552 vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_276_Right_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15038__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ net511 _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__or2_1
X_17976_ net639 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__inv_2
XANTENNA__19516__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14295__A2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19715_ clknet_leaf_35_clk game.writer.tracker.next_frame\[310\] net1340 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[310\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_29_Left_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16927_ _02359_ _02636_ net714 vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__o21a_1
XANTENNA__15980__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_291_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_358_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17233__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19646_ clknet_leaf_28_clk game.writer.tracker.next_frame\[241\] net1287 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[241\] sky130_fd_sc_hd__dfrtp_4
X_16858_ _02542_ net108 _02625_ net1725 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[243\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14596__B net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15809_ game.CPU.applesa.ab.check_walls.above.walls\[59\] net463 vssd1 vssd1 vccd1
+ vccd1 _01821_ sky130_fd_sc_hd__and2_1
XANTENNA__13255__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19577_ clknet_leaf_31_clk game.writer.tracker.next_frame\[172\] net1279 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[172\] sky130_fd_sc_hd__dfrtp_1
X_16789_ net146 _02466_ net105 _02598_ net2046 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[201\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__19666__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_338_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ net925 game.CPU.applesa.ab.absxs.body_x\[83\] game.CPU.applesa.ab.absxs.body_y\[80\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__a22o_1
XANTENNA__10608__A2 _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18528_ net601 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__inv_2
XANTENNA__11805__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09261_ game.CPU.randy.counter1.count\[5\] vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__inv_2
X_18459_ net654 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__inv_2
XANTENNA__11281__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16744__A1 _02299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Left_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_334_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_303_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15501__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Left_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_334_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13558__B2 game.writer.tracker.frame\[97\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09192_ game.CPU.applesa.ab.check_walls.above.walls\[115\] vssd1 vssd1 vccd1 vccd1
+ _03441_ sky130_fd_sc_hd__inv_2
XANTENNA_clkload60_A clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16316__B _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout219_A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_214_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10792__A1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15180__B1 _03197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1030_A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_302_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1128_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout490_A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16051__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout588_A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__A game.CPU.applesa.ab.check_walls.above.walls\[50\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold14 game.CPU.start_pause_button1.eD1.Q1 vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_328_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_243_Right_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19196__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08976_ game.CPU.applesa.ab.absxs.body_x\[5\] vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__inv_2
Xhold25 game.CPU.walls.abc.number\[1\] vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14286__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold36 game.CPU.kyle.L1.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_270_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold47 game.CPU.applesa.off_bc.Q1 vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11195__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold58 game.CPU.clock1.game_state\[1\] vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_279_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold69 net42 vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18259__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17224__A2 _02720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15599__A2_N net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16432__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11923__B net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout922_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16983__A1 _02461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09528_ net1157 game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1 vccd1
+ vccd1 _03771_ sky130_fd_sc_hd__or2_1
XANTENNA__15114__C net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12100__A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18990__Q game.CPU.applesa.ab.check_walls.above.walls\[35\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ net923 game.CPU.applesa.ab.absxs.body_x\[70\] game.CPU.applesa.ab.absxs.body_y\[69\]
+ net899 _03695_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__o221a_1
XANTENNA__16735__A1 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12470_ game.CPU.applesa.ab.absxs.body_x\[13\] net378 net366 game.CPU.applesa.ab.absxs.body_y\[15\]
+ _06340_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_314_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16226__B net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_340_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11421_ net798 net315 vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_152_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_340_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14140_ _07826_ _07831_ _07906_ _07938_ _07994_ vssd1 vssd1 vccd1 vccd1 _08014_ sky130_fd_sc_hd__o2111a_1
X_11352_ net773 _05240_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_278_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17160__A1 _02444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16513__Y _02455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10303_ _04482_ _04484_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__nand2_4
X_14071_ net961 game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 _07945_ sky130_fd_sc_hd__or2_1
X_11283_ _05171_ _05172_ _04930_ _05006_ _05169_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__o2111a_1
X_13022_ net484 net697 _06879_ _06895_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__a31o_1
XANTENNA__19539__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ game.CPU.applesa.ab.count_luck\[2\] game.CPU.applesa.ab.count_luck\[0\] _04425_
+ game.CPU.applesa.ab.count_luck\[1\] vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_91_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10535__A1 game.CPU.applesa.ab.absxs.body_x\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_258_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1001 net1009 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
Xfanout1012 net1013 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_4
X_17830_ _03150_ _03159_ _03160_ _03146_ net2051 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__a32o_1
XANTENNA__09127__Y _03376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10165_ net1078 _04359_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__or2_1
Xfanout1023 net1025 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_238_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1034 net1041 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_210_Right_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1045 net1051 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__buf_6
XFILLER_0_246_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1056 net1059 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_163_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17761_ _03116_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__inv_2
XANTENNA__13485__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1067 net1068 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__buf_4
X_14973_ net1226 net1253 game.CPU.applesa.ab.check_walls.above.walls\[1\] vssd1 vssd1
+ vccd1 vccd1 _00287_ sky130_fd_sc_hd__and3_1
XANTENNA__18563__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ _04301_ _04303_ _04266_ _04298_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__a211o_1
XANTENNA__19689__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__buf_4
X_19500_ clknet_leaf_25_clk game.writer.tracker.next_frame\[95\] net1319 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[95\] sky130_fd_sc_hd__dfrtp_1
Xfanout1089 net1090 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_4
X_16712_ net161 net69 net106 _02571_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[151\]
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17215__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13924_ _07793_ _07794_ _07789_ _07791_ vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__a211o_1
X_17692_ game.CPU.walls.rand_wall.count_luck\[6\] _03071_ net1856 vssd1 vssd1 vccd1
+ vccd1 _03073_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_214_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19431_ clknet_leaf_39_clk game.writer.tracker.next_frame\[26\] net1352 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_254_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16643_ net114 net157 _02539_ net727 vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__o31a_1
XANTENNA__11833__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13855_ net279 _07722_ _07723_ net484 vssd1 vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__a31o_1
XANTENNA__16974__A1 _02450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19061__Q game.CPU.applesa.ab.check_walls.above.walls\[106\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12806_ game.writer.tracker.frame\[330\] game.writer.tracker.frame\[331\] net998
+ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19362_ clknet_leaf_68_clk _01368_ _00943_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_16574_ net230 _02417_ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__nor2_4
XANTENNA__09303__B game.CPU.applesa.ab.absxs.body_x\[55\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13786_ net285 _07644_ _07650_ _07659_ net242 vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__a311o_1
XANTENNA__15024__C game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10998_ game.CPU.applesa.ab.absxs.body_x\[45\] net413 vssd1 vssd1 vccd1 vccd1 _04888_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_347_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11799__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10449__B net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18313_ net620 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__inv_2
X_15525_ _01524_ _01546_ _01506_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__a21o_1
XANTENNA__16726__A1 _02359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12737_ game.writer.tracker.frame\[72\] game.writer.tracker.frame\[73\] net1014 vssd1
+ vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_270_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_252_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19293_ clknet_leaf_71_clk _01337_ _00912_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.off_bc.D
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18244_ net645 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
XFILLER_0_270_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15456_ _01435_ _01440_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_174_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ game.CPU.luck1.Qa\[0\] net1274 _04733_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__mux2_1
XANTENNA__14201__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19069__CLK net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_316_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_316_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15040__B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14407_ game.CPU.applesa.ab.absxs.body_y\[44\] net986 vssd1 vssd1 vccd1 vccd1 _08281_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__11015__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ game.CPU.applesa.ab.check_walls.above.walls\[187\] net761 vssd1 vssd1 vccd1
+ vccd1 _05508_ sky130_fd_sc_hd__xnor2_2
X_18175_ net603 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__inv_2
XFILLER_0_288_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15387_ _08927_ _08928_ vssd1 vssd1 vccd1 vccd1 _08929_ sky130_fd_sc_hd__nor2_1
XANTENNA__10465__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_345_Right_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12599_ game.CPU.applesa.ab.absxs.body_y\[109\] net524 net378 game.CPU.applesa.ab.absxs.body_x\[109\]
+ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_142_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17126_ net156 _02382_ net76 _02710_ net1658 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[426\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14338_ game.CPU.applesa.ab.absxs.body_x\[39\] net873 net963 _03312_ vssd1 vssd1
+ vccd1 vccd1 _08212_ sky130_fd_sc_hd__o22a_1
XANTENNA__17151__A1 _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold506 game.writer.tracker.frame\[15\] vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_296_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16423__Y _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold517 game.CPU.applesa.twoapples.count_luck\[2\] vssd1 vssd1 vccd1 vccd1 net1902
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 game.writer.tracker.frame\[385\] vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_296_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17057_ _02428_ net84 _02687_ net1557 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[380\]
+ sky130_fd_sc_hd__a22o_1
Xhold539 game.writer.tracker.frame\[518\] vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14269_ game.CPU.applesa.ab.absxs.body_x\[48\] net889 net858 game.CPU.applesa.ab.absxs.body_y\[51\]
+ vssd1 vssd1 vccd1 vccd1 _08143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_284_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16008_ game.CPU.applesa.ab.absxs.body_y\[60\] net453 vssd1 vssd1 vccd1 vccd1 _02020_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_55_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_263_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12920__C1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__A1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18906__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__B2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14268__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ net648 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_302_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17206__A2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_224_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11743__B net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19629_ clknet_leaf_26_clk game.writer.tracker.next_frame\[224\] net1311 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[224\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16965__A1 _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15768__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout169_A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_274_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09313_ net1094 game.CPU.applesa.ab.absxs.body_x\[66\] vssd1 vssd1 vccd1 vccd1 _03556_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_46_Left_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11254__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16717__A1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_216_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16327__A _06573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout336_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13450__S net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_60_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_346_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_196_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09244_ game.CPU.applesa.twoapples.good_spot vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1078_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14256__A1_N net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09175_ game.CPU.applesa.ab.check_walls.above.walls\[81\] vssd1 vssd1 vccd1 vccd1
+ _03424_ sky130_fd_sc_hd__inv_2
XFILLER_0_334_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10375__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout124_X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout503_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_312_Right_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13951__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17142__A1 _02413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13951__B2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15885__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10765__B2 game.CPU.applesa.ab.absxs.body_y\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11962__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17158__A _02237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput15 net15 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Left_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput26 net1278 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
Xoutput37 net37 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_113_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_285_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout872_A _03374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__A1 _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18586__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10822__B game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_227_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19831__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16653__B1 _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18985__Q game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08959_ game.CPU.apple_location\[3\] vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__inv_2
XANTENNA__11934__A game.CPU.applesa.ab.check_walls.above.walls\[165\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11970_ _05426_ _05428_ _05429_ _05430_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__or4_1
XANTENNA__09686__A2 game.CPU.applesa.ab.absxs.body_y\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16405__B1 _02375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19981__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ net1166 _04367_ _04813_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__a21o_1
XANTENNA__16956__A1 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14527__B1_N _07742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_316_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Left_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_329_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13640_ game.writer.tracker.frame\[61\] game.writer.tracker.frame\[63\] game.writer.tracker.frame\[64\]
+ game.writer.tracker.frame\[62\] net980 net1040 vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__mux4_1
XANTENNA__16420__A3 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10852_ _04750_ _04751_ _04754_ _04741_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__a31o_1
XFILLER_0_329_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_296_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16508__Y _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14431__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12978__C1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_238_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13571_ _07441_ _07444_ net203 vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__mux2_1
X_10783_ _03308_ net327 vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__nor2_1
XANTENNA__11245__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13360__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_344_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_325_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15141__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15310_ game.CPU.applesa.twomode.number\[7\] _08851_ net757 vssd1 vssd1 vccd1 vccd1
+ _08857_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ game.CPU.applesa.ab.absxs.body_y\[70\] net522 vssd1 vssd1 vccd1 vccd1 _06399_
+ sky130_fd_sc_hd__xnor2_1
X_16290_ _02274_ _02291_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__or2_1
XANTENNA__16184__A2 _02190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15241_ game.CPU.kyle.L1.cnt_500hz\[3\] _08801_ vssd1 vssd1 vccd1 vccd1 _08802_ sky130_fd_sc_hd__and2_1
X_12453_ game.CPU.applesa.ab.absxs.body_y\[51\] net367 vssd1 vssd1 vccd1 vccd1 _06330_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_313_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_313_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19361__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ game.CPU.applesa.ab.check_walls.above.walls\[95\] net260 net316 net806 vssd1
+ vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_124_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15172_ game.CPU.bodymain1.main.score\[7\] game.CPU.bodymain1.main.score\[5\] vssd1
+ vssd1 vccd1 vccd1 _08748_ sky130_fd_sc_hd__and2b_1
X_12384_ _03353_ net369 vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__nor2_1
XANTENNA__17133__A1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_340_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Left_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17068__A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14123_ net1058 _03392_ _03395_ net945 _07996_ vssd1 vssd1 vccd1 vccd1 _07997_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11335_ _05223_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__inv_2
XANTENNA__18929__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_327_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19980_ clknet_leaf_42_clk game.writer.tracker.next_frame\[575\] net1326 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[575\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_266_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14498__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_265_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18931_ clknet_leaf_4_clk net1399 _00615_ vssd1 vssd1 vccd1 vccd1 game.CPU.start_pause_button1.eD1.Q2
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_249_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14054_ net983 net790 vssd1 vssd1 vccd1 vccd1 _07928_ sky130_fd_sc_hd__nand2_1
X_11266_ game.CPU.applesa.ab.absxs.body_x\[100\] net415 net397 game.CPU.applesa.ab.absxs.body_y\[103\]
+ _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__a221o_1
XANTENNA__17510__A_N _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13005_ game.writer.tracker.frame\[572\] game.writer.tracker.frame\[573\] net1021
+ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__mux2_1
X_10217_ _04392_ _04399_ _04393_ _04389_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__o211a_1
XFILLER_0_281_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18862_ clknet_leaf_1_clk _01253_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_11197_ game.CPU.applesa.ab.absxs.body_x\[20\] net415 vssd1 vssd1 vccd1 vccd1 _05087_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_246_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17813_ _01438_ _01444_ _08897_ _08936_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13458__A0 _06985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10148_ net1260 game.CPU.randy.f1.state\[4\] vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__nand2b_1
X_18793_ clknet_leaf_4_clk _01208_ _00530_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[5\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_265_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15998__A2 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11844__A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13553__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17744_ _03100_ game.CPU.applesa.ab.count\[3\] game.CPU.applesa.ab.count\[1\] game.CPU.applesa.ab.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__and4b_1
X_10079_ _04225_ _04270_ _04228_ _04215_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o211a_1
X_14956_ _08729_ _08732_ _08731_ _08724_ vssd1 vssd1 vccd1 vccd1 _08733_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_50_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Left_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09314__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ net1044 game.CPU.applesa.ab.check_walls.above.walls\[123\] vssd1 vssd1 vccd1
+ vccd1 _07781_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17675_ _03523_ _03060_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__nor2_1
XANTENNA__15035__B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_338_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16947__A1 _02391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14887_ net1125 _08430_ vssd1 vssd1 vccd1 vccd1 _08664_ sky130_fd_sc_hd__nor2_1
XFILLER_0_348_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19414_ clknet_leaf_47_clk game.writer.tracker.next_frame\[9\] net1295 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[9\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11758__A2_N net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16626_ net113 _02531_ net714 vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__o21a_1
XANTENNA__13305__S0 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13838_ game.writer.tracker.frame\[517\] game.writer.tracker.frame\[519\] game.writer.tracker.frame\[520\]
+ game.writer.tracker.frame\[518\] net971 net1008 vssd1 vssd1 vccd1 vccd1 _07712_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__16411__A3 _02379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14422__A2 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_308_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19345_ clknet_leaf_72_clk _01360_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.count\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16557_ net1945 _02481_ _02485_ net125 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[82\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12433__A1 game.CPU.applesa.ab.absxs.body_y\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13769_ net498 _07641_ _07642_ vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__and3_1
XANTENNA__12675__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12433__B2 game.CPU.applesa.ab.absxs.body_y\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_42_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_186_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15051__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15508_ net888 net1057 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12984__A2 _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19276_ clknet_leaf_7_clk _00046_ _00906_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_16488_ net2055 _02433_ _02435_ _02273_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[63\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19704__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18227_ net664 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15439_ _08914_ _08927_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__or2_1
XANTENNA__14186__B2 game.CPU.applesa.ab.absxs.body_x\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14890__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_300_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13933__A1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18158_ net630 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__inv_2
XANTENNA__13933__B2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17124__A1 _02378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_349_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold303 game.writer.tracker.frame\[566\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_211_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17109_ _02577_ net81 _02705_ net1830 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[414\]
+ sky130_fd_sc_hd__a22o_1
Xhold314 game.writer.tracker.frame\[163\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 game.writer.tracker.frame\[217\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19854__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18089_ net605 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__inv_2
XANTENNA__10482__X _04609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold336 game.writer.tracker.frame\[471\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_257_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 game.CPU.walls.rand_wall.count1 vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold358 game.writer.tracker.frame\[565\] vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_269_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold369 game.CPU.randy.counter1.count\[4\] vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ net1109 net1262 vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__nand2_1
XANTENNA__11738__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout805 game.CPU.applesa.ab.check_walls.above.walls\[94\] vssd1 vssd1 vccd1 vccd1
+ net805 sky130_fd_sc_hd__clkbuf_4
Xfanout816 game.CPU.applesa.ab.check_walls.above.walls\[63\] vssd1 vssd1 vccd1 vccd1
+ net816 sky130_fd_sc_hd__buf_4
X_20051_ net1369 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
X_09862_ net1103 game.CPU.applesa.ab.absxs.body_x\[45\] vssd1 vssd1 vccd1 vccd1 _04105_
+ sky130_fd_sc_hd__xor2_1
Xfanout827 game.CPU.applesa.ab.check_walls.above.walls\[23\] vssd1 vssd1 vccd1 vccd1
+ net827 sky130_fd_sc_hd__buf_2
XFILLER_0_309_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout838 net839 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16610__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_271_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout849 _04157_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__buf_2
XFILLER_0_252_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09793_ net1143 game.CPU.applesa.ab.absxs.body_y\[42\] vssd1 vssd1 vccd1 vccd1 _04036_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout286_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16650__A3 _02412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14130__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_222_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09224__A game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11473__B net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16938__A1 _02375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout453_A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1195_A game.CPU.walls.rand_wall.good_spot vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_327_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13847__S1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_326_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout241_X net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12585__A game.CPU.applesa.ab.absxs.body_y\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_341_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_33_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19384__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14177__B2 game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09227_ game.CPU.applesa.ab.check_walls.above.walls\[178\] vssd1 vssd1 vccd1 vccd1
+ _03476_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_311_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1150_X net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_307_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1248_X net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09158_ game.CPU.applesa.ab.check_walls.above.walls\[50\] vssd1 vssd1 vccd1 vccd1
+ _03407_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17159__Y _02720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_233_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10738__B2 game.CPU.applesa.ab.absxs.body_y\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16504__B _02400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09089_ game.CPU.applesa.ab.absxs.body_y\[58\] vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14305__A game.CPU.applesa.ab.absxs.body_x\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09570__A2_N game.CPU.applesa.ab.absxs.body_x\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11120_ _03282_ net544 vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__nand2_1
XANTENNA__16874__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11648__B net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09356__A1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11051_ _03253_ net320 vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09356__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16626__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ net1165 game.CPU.applesa.out_random_2\[1\] vssd1 vssd1 vccd1 vccd1 _04210_
+ sky130_fd_sc_hd__nand2_2
XANTENNA__10271__C game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_322_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _08619_ _08620_ net138 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__and3b_1
XANTENNA__15136__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11664__A game.CPU.applesa.ab.check_walls.above.walls\[120\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14101__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14101__B2 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15790_ game.CPU.applesa.ab.absxs.body_x\[72\] net356 vssd1 vssd1 vccd1 vccd1 _01802_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_270_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12479__B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09134__A game.CPU.applesa.ab.check_walls.above.walls\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14741_ _08567_ _08568_ net55 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__and3b_1
XANTENNA__16929__A1 _02512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11953_ net569 _05301_ _05836_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__and3_1
XANTENNA__13860__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16929__B2 game.writer.tracker.frame\[289\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18447__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10904_ game.CPU.applesa.ab.check_walls.collision_down _04799_ _04801_ game.CPU.applesa.ab.check_walls.collision_right
+ _04805_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_86_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17351__A _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17460_ _04638_ _02784_ _02798_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__and3_1
XANTENNA__18601__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14672_ _08510_ _08507_ _08506_ vssd1 vssd1 vccd1 vccd1 _08511_ sky130_fd_sc_hd__or3b_1
XANTENNA__19727__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11884_ net827 net312 vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__or2_1
XFILLER_0_345_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13838__S1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16411_ net135 net115 _02379_ net556 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a31oi_2
XTAP_TAPCELL_ROW_28_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13623_ game.writer.tracker.frame\[277\] game.writer.tracker.frame\[279\] game.writer.tracker.frame\[280\]
+ game.writer.tracker.frame\[278\] net976 net1018 vssd1 vssd1 vccd1 vccd1 _07497_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835_ game.CPU.speed1.Qa\[0\] game.CPU.speed1.Qa\[2\] _04736_ vssd1 vssd1 vccd1
+ vccd1 _00014_ sky130_fd_sc_hd__mux2_1
X_17391_ _02783_ _02820_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_24_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_251_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19130_ net1184 _00171_ _00801_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[175\]
+ sky130_fd_sc_hd__dfrtp_4
X_16342_ _02279_ _02295_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__nand2_2
X_13554_ game.writer.tracker.frame\[65\] game.writer.tracker.frame\[67\] game.writer.tracker.frame\[68\]
+ game.writer.tracker.frame\[66\] net978 net1026 vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_158_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10766_ game.CPU.applesa.ab.absxs.body_y\[82\] _04673_ _04674_ game.CPU.applesa.ab.absxs.body_y\[78\]
+ vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_333_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10727__B _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_332_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12411__A2_N net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19061_ net1190 _00095_ _00732_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[106\]
+ sky130_fd_sc_hd__dfrtp_4
X_12505_ game.CPU.applesa.ab.absxs.body_x\[74\] net374 vssd1 vssd1 vccd1 vccd1 _06382_
+ sky130_fd_sc_hd__xnor2_1
X_16273_ net2044 _02260_ _02267_ _02273_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[5\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18751__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19877__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13485_ net477 _07109_ net693 vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__a21o_1
X_10697_ game.CPU.applesa.ab.absxs.body_y\[85\] _04610_ _04611_ game.CPU.applesa.ab.absxs.body_y\[81\]
+ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__a22o_1
XANTENNA__12179__B1 _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18012_ net648 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__inv_2
X_15224_ game.CPU.applesa.normal1.number\[5\] _08783_ vssd1 vssd1 vccd1 vccd1 _08789_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__17069__Y _02693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13597__Y _07471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12436_ _03253_ net372 vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17106__A1 _02576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10729__A1 game.CPU.applesa.ab.absxs.body_y\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_124_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16414__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10729__B2 game.CPU.applesa.ab.absxs.body_y\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13391__A2 _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15155_ net1214 net1239 net783 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__and3_1
X_12367_ _06234_ _06235_ _06240_ _06243_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_97_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14106_ net1073 game.CPU.applesa.ab.check_walls.above.walls\[48\] vssd1 vssd1 vccd1
+ vccd1 _07980_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_266_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11318_ _05194_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__nor2_4
X_19963_ clknet_leaf_43_clk game.writer.tracker.next_frame\[558\] net1306 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[558\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_266_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15086_ net1206 net1232 game.CPU.applesa.ab.check_walls.above.walls\[114\] vssd1
+ vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__and3_1
X_12298_ net827 net421 vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__or2_1
XFILLER_0_276_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14037_ net882 game.CPU.applesa.ab.check_walls.above.walls\[113\] net796 net856 vssd1
+ vssd1 vccd1 vccd1 _07911_ sky130_fd_sc_hd__o22a_1
X_18914_ clknet_leaf_5_clk net1395 _00598_ vssd1 vssd1 vccd1 vccd1 game.CPU.up_button.eD1.Q1
+ sky130_fd_sc_hd__dfrtp_1
X_11249_ game.CPU.applesa.ab.absxs.body_y\[7\] net397 vssd1 vssd1 vccd1 vccd1 _05139_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_253_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16880__A3 _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19894_ clknet_leaf_14_clk game.writer.tracker.next_frame\[489\] net1283 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[489\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09898__A2 _03825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16617__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_182_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18845_ clknet_leaf_0_clk _01236_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11574__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18776_ clknet_leaf_69_clk _01193_ _00513_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[86\]
+ sky130_fd_sc_hd__dfrtp_4
X_15988_ _03419_ net447 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12389__B net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17727_ game.CPU.applesa.ab.count_luck\[5\] _03093_ _03085_ vssd1 vssd1 vccd1 vccd1
+ _03095_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09044__A game.CPU.applesa.ab.absxs.body_y\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14939_ _08680_ _08682_ vssd1 vssd1 vccd1 vccd1 _08716_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13851__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_340_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17042__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17658_ game.CPU.kyle.L1.cnt_500hz\[9\] _03047_ game.CPU.kyle.L1.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__a21o_1
XFILLER_0_348_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16609_ net1518 _02515_ _02519_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[99\]
+ sky130_fd_sc_hd__a21o_1
X_17589_ net1478 _03009_ net582 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_63_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_271_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_15_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_308_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19328_ clknet_leaf_72_clk net1428 _00933_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twomode.number\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_193_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14159__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14159__B2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19259_ clknet_leaf_57_clk _01327_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.count_luck\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16605__A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18092__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_311_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09012_ game.CPU.applesa.ab.absxs.body_x\[97\] vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13948__B game.CPU.applesa.ab.check_walls.above.walls\[135\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15936__A2_N net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11917__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold100 game.CPU.walls.rand_wall.count\[1\] vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold111 game.writer.tracker.frame\[310\] vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold122 game.writer.tracker.frame\[373\] vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 game.writer.tracker.frame\[99\] vssd1 vssd1 vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 game.writer.tracker.frame\[437\] vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16856__B1 _02623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_269_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12590__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09219__A game.CPU.applesa.ab.check_walls.above.walls\[165\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 game.writer.tracker.frame\[167\] vssd1 vssd1 vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 game.CPU.randy.f1.c1.count\[16\] vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 game.writer.tracker.frame\[170\] vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_282_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold188 game.writer.tracker.frame\[207\] vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 game.writer.tracker.frame\[205\] vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 net604 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_4
X_09914_ net1263 game.CPU.bodymain1.main.pause_clk vssd1 vssd1 vccd1 vccd1 _04156_
+ sky130_fd_sc_hd__and2_4
Xfanout613 net614 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_4
XANTENNA__16871__A3 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_272_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout624 net625 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1110_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout635 net636 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_298_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1208_A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20034_ net1382 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_95_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout646 net651 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_2
Xfanout657 net658 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__buf_4
X_09845_ _04086_ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__nand2_1
XANTENNA_input6_A gpio_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout191_X net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 net670 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__buf_4
Xfanout679 net680 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout668_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14095__B1 _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18624__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ net906 net1172 net1170 net902 _04018_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__a221o_4
XANTENNA__16994__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12299__B _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13842__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18267__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1198_X net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12586__Y _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_293_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18774__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_235_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10620_ _04174_ _04176_ _04581_ _04606_ net328 vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a41o_4
XFILLER_0_76_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15122__C game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10551_ _03279_ net330 vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13270_ game.writer.tracker.frame\[496\] game.writer.tracker.frame\[497\] net998
+ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__mux2_1
X_10482_ net849 _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout992_X net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16234__B _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_322_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11659__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12221_ _06103_ _06104_ _06105_ _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__or4_1
XANTENNA__10563__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14035__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14570__B2 game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__B2 game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09129__A game.CPU.applesa.ab.check_walls.above.walls\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12152_ _06036_ _06037_ _06038_ _06035_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__a211o_1
XANTENNA__11378__B net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_248_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11103_ _03216_ net404 vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09329__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13874__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16960_ _02419_ net94 net559 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_246_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17346__A _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12083_ game.CPU.applesa.ab.check_walls.above.walls\[20\] net555 vssd1 vssd1 vccd1
+ vccd1 _05970_ sky130_fd_sc_hd__nand2_1
XANTENNA__16250__A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_263_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11034_ game.CPU.applesa.ab.absxs.body_y\[67\] net399 vssd1 vssd1 vccd1 vccd1 _04924_
+ sky130_fd_sc_hd__xnor2_1
X_15911_ game.CPU.applesa.ab.check_walls.above.walls\[128\] net269 vssd1 vssd1 vccd1
+ vccd1 _01923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_263_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16891_ _02460_ net93 _02639_ net1564 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[262\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_235_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_188_Right_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17272__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18630_ clknet_leaf_10_clk _01047_ _00367_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09135__Y _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15842_ game.CPU.applesa.ab.check_walls.above.walls\[20\] net453 vssd1 vssd1 vccd1
+ vccd1 _01854_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_246_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18561_ clknet_leaf_8_clk _00981_ _00298_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_15773_ game.CPU.applesa.ab.absxs.body_y\[104\] net452 vssd1 vssd1 vccd1 vccd1 _01785_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12985_ _06822_ _06858_ _06703_ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12002__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13813__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17512_ _02916_ _02917_ _02918_ _02940_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__a31o_1
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14724_ game.CPU.randy.counter1.count1\[7\] _08555_ vssd1 vssd1 vccd1 vccd1 _08557_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_335_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ net748 _05587_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__nand2_1
X_18492_ net617 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_358_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17443_ game.CPU.kyle.L1.nextState\[5\] game.CPU.kyle.L1.nextState\[4\] _02827_ vssd1
+ vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__nand3_4
XFILLER_0_156_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14655_ net753 _08489_ _08491_ vssd1 vssd1 vccd1 vccd1 _08494_ sky130_fd_sc_hd__and3b_1
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11867_ net751 _05397_ _05399_ net574 vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ game.writer.tracker.frame\[289\] game.writer.tracker.frame\[291\] game.writer.tracker.frame\[292\]
+ game.writer.tracker.frame\[290\] net967 net996 vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__mux4_1
XFILLER_0_184_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17374_ _02793_ _02797_ _02803_ _02795_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a22o_1
X_10818_ game.CPU.applesa.ab.absxs.body_y\[11\] _04689_ _04707_ game.CPU.applesa.ab.absxs.body_y\[7\]
+ vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__a22o_1
XANTENNA__15032__C net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14586_ game.CPU.clock1.counter\[5\] game.CPU.clock1.counter\[8\] vssd1 vssd1 vccd1
+ vccd1 _08448_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ game.CPU.applesa.ab.check_walls.above.walls\[196\] net392 _05684_ _05685_
+ _05443_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a2111o_1
X_19113_ net1181 _00152_ _00784_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[158\]
+ sky130_fd_sc_hd__dfrtp_4
X_16325_ net70 _02318_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__nor2_1
X_13537_ game.writer.tracker.frame\[81\] game.writer.tracker.frame\[83\] game.writer.tracker.frame\[84\]
+ game.writer.tracker.frame\[82\] net978 net1028 vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_99_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10749_ game.CPU.applesa.ab.absxs.body_y\[114\] _04663_ _04664_ game.CPU.applesa.ab.absxs.body_y\[110\]
+ vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__a22o_1
X_19044_ net1191 _00275_ _00715_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[89\]
+ sky130_fd_sc_hd__dfrtp_4
X_16256_ net1008 _08400_ _02261_ net865 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__o211a_1
X_13468_ net495 _07079_ net684 vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15207_ game.CPU.applesa.normal1.number\[6\] _08770_ vssd1 vssd1 vccd1 vccd1 _08775_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09568__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ game.CPU.applesa.ab.absxs.body_x\[35\] net528 net518 game.CPU.applesa.ab.absxs.body_y\[34\]
+ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09568__B2 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10473__A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16187_ _01681_ _01682_ _01683_ _02198_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_346_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13399_ _06874_ _06890_ net685 vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15138_ net1210 net1236 net787 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__and3_1
XANTENNA__15983__B net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13784__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13747__S0 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19946_ clknet_leaf_33_clk game.writer.tracker.next_frame\[541\] net1324 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[541\] sky130_fd_sc_hd__dfrtp_1
X_15069_ net1217 net1246 game.CPU.applesa.ab.check_walls.above.walls\[97\] vssd1 vssd1
+ vccd1 vccd1 _00094_ sky130_fd_sc_hd__and3_1
XFILLER_0_294_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__18647__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Left_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19877_ clknet_leaf_27_clk game.writer.tracker.next_frame\[472\] net1316 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[472\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10886__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ net1100 _03283_ game.CPU.applesa.ab.absxs.body_y\[16\] net895 _03871_ vssd1
+ vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__a221o_1
X_18828_ clknet_leaf_1_clk _01219_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.lcd_rs
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__14077__B1 game.CPU.applesa.ab.YMAX\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09561_ net1161 game.CPU.applesa.ab.absxs.body_y\[60\] vssd1 vssd1 vccd1 vccd1 _03804_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__13824__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18759_ clknet_leaf_12_clk _01176_ _00496_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[53\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__18087__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_357_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09492_ net1097 _03480_ _03482_ net1145 _03730_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__a221o_1
XFILLER_0_222_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout151_A _02270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10648__A game.CPU.bad_collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16606__Y _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_351_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13959__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16335__A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1060_A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1158_A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_320_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12582__B net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19422__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_230_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11479__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13879__A1_N net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout204_X net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1325_A net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11198__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15893__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_A game.CPU.applesa.ab.check_walls.above.walls\[172\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13694__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13738__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1113_X net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12315__B1 _06122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout410 net411 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_4
XANTENNA__19572__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout421 _04782_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_245_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout432 net437 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_8
Xfanout443 _08429_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_4
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_6
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout952_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 net470 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_4
XANTENNA__14302__B net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16057__A1 net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout476 net480 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09731__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16057__B2 net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20017_ net1277 vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
Xfanout487 net489 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_4
X_09828_ net1102 game.CPU.applesa.ab.absxs.body_x\[13\] vssd1 vssd1 vccd1 vccd1 _04071_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__09731__B2 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout498 net499 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout64_A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10341__A2 _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_241_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09759_ net1103 game.CPU.applesa.ab.check_walls.above.walls\[25\] vssd1 vssd1 vccd1
+ vccd1 _04002_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_240_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16114__A1_N net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12770_ game.writer.tracker.frame\[88\] game.writer.tracker.frame\[89\] net1028 vssd1
+ vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__mux2_1
XANTENNA__12443__A1_N game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17557__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16229__B net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ net813 net307 net304 net812 vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__a22o_1
XANTENNA__15133__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11841__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ game.CPU.applesa.ab.absxs.body_x\[90\] net1053 vssd1 vssd1 vccd1 vccd1 _08314_
+ sky130_fd_sc_hd__or2_1
X_11652_ net744 _05538_ _05540_ net567 vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__a22o_1
XANTENNA__16780__A2 _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17309__B2 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout61 net65 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_2
Xfanout72 _02691_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_4
X_10603_ game.CPU.applesa.ab.absxs.body_x\[90\] _04590_ net329 game.CPU.applesa.ab.absxs.body_x\[86\]
+ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout83 net84 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_2
X_14371_ _08241_ _08242_ _08243_ _08244_ vssd1 vssd1 vccd1 vccd1 _08245_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_155_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout94 net96 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_2
X_11583_ _05423_ _05439_ _05453_ _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_330_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_308_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire833 _08938_ vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_1
X_16110_ game.CPU.applesa.ab.check_walls.above.walls\[11\] net462 net447 game.CPU.applesa.ab.check_walls.above.walls\[13\]
+ _01689_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__o221a_1
X_13322_ net493 _06720_ _07195_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__a21o_1
X_17090_ _02322_ _02693_ net737 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__o21a_1
X_10534_ net754 _04639_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_21_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12492__B net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16041_ _03311_ net453 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__nand2_1
XFILLER_0_311_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13253_ _07122_ _07123_ _07125_ _07124_ net487 net683 vssd1 vssd1 vccd1 vccd1 _07127_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_257_Right_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10465_ net1266 _04595_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__and2_1
XFILLER_0_161_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16532__X _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12554__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12204_ _05944_ _06088_ _06089_ _05945_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__or4b_1
XANTENNA__19915__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13184_ net231 _07057_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_94_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10396_ _04350_ _04353_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__nor2_1
XFILLER_0_310_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19800_ clknet_leaf_33_clk game.writer.tracker.next_frame\[395\] net1324 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[395\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11676__X _05565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10580__X _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12135_ _03418_ net553 vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__xnor2_1
X_17992_ net640 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__inv_2
XANTENNA__13503__C1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19731_ clknet_leaf_19_clk game.writer.tracker.next_frame\[326\] net1337 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[326\] sky130_fd_sc_hd__dfrtp_1
X_16943_ _02379_ net87 net556 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11836__B net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ net795 net386 vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_166_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10740__B _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_341_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14212__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11017_ _04903_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__or2_2
X_16874_ net157 _02432_ net99 net729 vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__o31a_1
X_19662_ clknet_leaf_23_clk game.writer.tracker.next_frame\[257\] net1344 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[257\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09306__B game.CPU.applesa.ab.absxs.body_x\[54\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15027__C net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15825_ game.CPU.applesa.ab.absxs.body_x\[89\] net471 net431 game.CPU.applesa.ab.absxs.body_y\[91\]
+ _01836_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__o221a_1
X_18613_ clknet_leaf_70_clk _01030_ _00350_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[99\]
+ sky130_fd_sc_hd__dfrtp_4
X_19593_ clknet_leaf_37_clk game.writer.tracker.next_frame\[188\] net1355 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[188\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17260__A3 _02619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12609__B2 game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18544_ net611 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__inv_2
X_15756_ game.CPU.applesa.ab.absxs.body_x\[20\] net356 vssd1 vssd1 vccd1 vccd1 _01768_
+ sky130_fd_sc_hd__xnor2_1
X_12968_ _06654_ _06657_ net682 vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_231_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12667__B _06487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ _03517_ net54 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__and2_1
XANTENNA__11571__B net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15043__B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ game.CPU.applesa.ab.check_walls.above.walls\[14\] net302 _05805_ _05806_
+ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__a211o_1
X_18475_ net638 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11832__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15687_ _03226_ net356 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__nand2_1
X_12899_ _06771_ _06772_ net513 vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__mux2_1
X_17426_ _02779_ _02828_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14638_ _08480_ _08481_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[18\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15978__B net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16771__A2 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_177_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13585__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19445__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17357_ _02771_ _02776_ _02785_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14569_ net929 net1264 vssd1 vssd1 vccd1 vccd1 _08433_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_190_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_303_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16308_ _06572_ net835 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__nor2_1
X_17288_ net130 _02579_ net722 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__o21a_1
XFILLER_0_302_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload20 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__inv_16
XFILLER_0_70_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19027_ net1193 _00257_ _00698_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[72\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16239_ net967 _02245_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__nand2_1
Xclkload31 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload31/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload42 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__inv_6
XFILLER_0_341_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_224_Right_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload53 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload53/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__16442__X _02403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload64 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__inv_12
XANTENNA__19595__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09410__B1 game.CPU.applesa.ab.check_walls.above.walls\[135\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_266_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08992_ game.CPU.applesa.ab.absxs.body_x\[52\] vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_208_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10931__A game.CPU.applesa.ab.absxs.body_x\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_282_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13196__S1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19929_ clknet_leaf_48_clk game.writer.tracker.next_frame\[524\] net1302 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[524\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17236__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_305_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_317_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09613_ _03849_ _03851_ _03852_ _03853_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__or4_1
XANTENNA__15798__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13453__S net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19351__D game.CPU.applesa.twoapples.absxs.next_head\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09544_ net919 net1172 _03785_ _03786_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__a22o_1
XANTENNA__13273__A1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17539__A1 net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_203_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_277_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16049__B net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09475_ net1137 _03479_ net783 net907 _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout533_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10378__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_290_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_219_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15888__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14222__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16762__A2 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16336__Y _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11036__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout700_A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout321_X net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__clkinv_8
XANTENNA_fanout1063_X net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18812__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18280__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ _03493_ net747 vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__nor2_1
XFILLER_0_277_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18988__Q game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_320_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13628__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _04368_ _04373_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_358_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1205 net1206 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10562__A2 _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_243_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1216 game.CPU.walls.rand_wall.start_enable vssd1 vssd1 vccd1 vccd1 net1216
+ sky130_fd_sc_hd__buf_4
XANTENNA__09407__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11656__B net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1227 net1228 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__buf_2
Xfanout240 net243 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_4
XANTENNA_fanout955_X net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1238 net1242 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__clkbuf_2
Xfanout251 _05210_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_4
Xfanout1249 net1257 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__buf_2
Xfanout262 _05195_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_260_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13940_ net944 game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1 vccd1
+ vccd1 _07814_ sky130_fd_sc_hd__xor2_1
Xfanout273 game.CPU.walls.rand_wall.abduyd.next_wall\[0\] vssd1 vssd1 vccd1 vccd1
+ net273 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_227_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout284 net287 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_4
XANTENNA__19318__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout67_X net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout295 _05858_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_4
X_13871_ _03371_ net1052 _07743_ _07744_ net1043 vssd1 vssd1 vccd1 vccd1 _07745_ sky130_fd_sc_hd__o221a_4
XTAP_TAPCELL_ROW_31_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11672__A game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15610_ _03346_ net444 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_319_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16450__B2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12822_ game.writer.tracker.frame\[356\] game.writer.tracker.frame\[357\] net1001
+ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__mux2_1
XANTENNA__15144__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16590_ _02430_ net144 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__nor2_2
XANTENNA__13264__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09142__A game.CPU.applesa.ab.check_walls.above.walls\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15541_ net943 net955 net699 _01547_ _01561_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__a311o_1
XANTENNA__11275__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19468__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12753_ game.writer.tracker.frame\[112\] game.writer.tracker.frame\[113\] net997
+ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__mux2_2
XFILLER_0_201_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14983__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_326_Right_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16202__A1 game.CPU.applesa.ab.check_walls.above.walls\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16202__B2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11704_ game.CPU.applesa.ab.check_walls.above.walls\[164\] net250 net314 game.CPU.applesa.ab.check_walls.above.walls\[165\]
+ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__o22a_1
X_18260_ net648 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
X_15472_ _01454_ _01498_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_194_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12684_ net943 _06556_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_328_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16753__A2 _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17211_ net146 _02375_ net75 _02733_ net1657 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[488\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__16246__Y _02254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14423_ _03259_ net1067 net871 game.CPU.applesa.ab.absxs.body_y\[108\] _08295_ vssd1
+ vssd1 vccd1 vccd1 _08297_ sky130_fd_sc_hd__o221a_1
XFILLER_0_355_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11635_ game.CPU.applesa.ab.check_walls.above.walls\[154\] net766 vssd1 vssd1 vccd1
+ vccd1 _05524_ sky130_fd_sc_hd__xnor2_2
X_18191_ net608 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__inv_2
XFILLER_0_343_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17142_ _02413_ _02693_ net736 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14354_ _03277_ net1070 net984 _03347_ _08226_ vssd1 vssd1 vccd1 vccd1 _08228_ sky130_fd_sc_hd__o221a_1
X_11566_ net792 net314 vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11404__A2_N net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16505__A2 _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17702__A1 game.CPU.walls.rand_wall.input2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13319__A2 _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13305_ game.writer.tracker.frame\[4\] game.writer.tracker.frame\[6\] game.writer.tracker.frame\[7\]
+ game.writer.tracker.frame\[5\] net969 net1002 vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17073_ _02267_ net59 _02694_ game.writer.tracker.frame\[389\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[389\] sky130_fd_sc_hd__a22o_1
X_10517_ _04358_ _04631_ net562 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__o21ai_4
X_14285_ game.CPU.applesa.ab.absxs.body_x\[85\] net881 net1044 _03231_ vssd1 vssd1
+ vccd1 vccd1 _08159_ sky130_fd_sc_hd__o22a_1
XFILLER_0_268_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11497_ game.CPU.applesa.ab.check_walls.above.walls\[170\] net766 vssd1 vssd1 vccd1
+ vccd1 _05386_ sky130_fd_sc_hd__xor2_1
XANTENNA__12008__A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16024_ game.CPU.applesa.ab.absxs.body_y\[92\] net451 vssd1 vssd1 vccd1 vccd1 _02036_
+ sky130_fd_sc_hd__xnor2_1
X_13236_ game.writer.tracker.frame\[476\] game.writer.tracker.frame\[477\] net1013
+ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__mux2_1
X_10448_ net1118 net1120 vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_343_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_311_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13538__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11847__A game.CPU.applesa.ab.check_walls.above.walls\[53\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13167_ net496 _07040_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__or2_1
XFILLER_0_268_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10379_ net914 game.CPU.apple_location2\[1\] _04530_ _04531_ net1263 vssd1 vssd1
+ vccd1 vccd1 _04532_ sky130_fd_sc_hd__o221a_1
XANTENNA__14223__A game.CPU.applesa.ab.absxs.body_x\[40\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_236_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09317__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12118_ _05381_ _05384_ _05386_ _05388_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__or4b_1
XANTENNA__13178__S1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11566__B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15038__B net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13098_ _06934_ _06936_ net687 vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17975_ net643 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19714_ clknet_leaf_36_clk game.writer.tracker.next_frame\[309\] net1340 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[309\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_284_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15606__X _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16926_ _02434_ _02643_ _02649_ net1835 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[287\]
+ sky130_fd_sc_hd__a22o_1
X_12049_ net817 net553 vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_251_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11502__A1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_284_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19645_ clknet_leaf_15_clk game.writer.tracker.next_frame\[240\] net1289 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[240\] sky130_fd_sc_hd__dfrtp_1
X_16857_ net158 _02539_ net99 net730 vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__o31a_1
XANTENNA__17233__A3 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16441__B2 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_253_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13126__X _07000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15054__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15808_ game.CPU.applesa.ab.check_walls.above.walls\[59\] net463 vssd1 vssd1 vccd1
+ vccd1 _01820_ sky130_fd_sc_hd__nor2_1
XANTENNA__13255__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16788_ net156 _02291_ net100 net727 vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__o31a_1
X_19576_ clknet_leaf_31_clk game.writer.tracker.next_frame\[171\] net1279 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[171\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09459__B1 game.CPU.applesa.ab.absxs.body_y\[69\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_354_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16992__A2 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12397__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09052__A game.CPU.applesa.ab.absxs.body_y\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15739_ _03473_ net332 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__xnor2_1
X_18527_ net601 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__inv_2
XANTENNA__11266__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14893__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_303_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09260_ game.CPU.randy.counter1.count1\[6\] vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__inv_2
X_18458_ net654 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14204__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13558__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09191_ game.CPU.applesa.ab.check_walls.above.walls\[114\] vssd1 vssd1 vccd1 vccd1
+ _03440_ sky130_fd_sc_hd__inv_2
X_17409_ game.CPU.kyle.L1.nextState\[5\] game.CPU.kyle.L1.nextState\[4\] game.CPU.kyle.L1.nextState\[3\]
+ game.CPU.kyle.L1.nextState\[2\] vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__and4b_1
XANTENNA__15501__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18389_ net618 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10926__A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload53_A clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_299_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_214_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18985__CLK net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout114_A _02243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10792__A2 game.CPU.applesa.ab.absxs.body_y\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13730__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14133__A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1023_A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11741__A1 _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09227__A game.CPU.applesa.ab.check_walls.above.walls\[178\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__B net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ game.CPU.applesa.ab.absxs.body_x\[6\] vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout483_A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 game.CPU.walls.abc.number\[2\] vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_102_Left_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold26 game.CPU.right_button.sync1.Q vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold37 game.CPU.applesa.normal1.number\[0\] vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold48 game.CPU.randy.f1.c1.count\[18\] vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 game.CPU.applesa.ab.absxs.body_x\[1\] vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_279_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout650_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout271_X net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19610__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16432__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16983__A2 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09527_ net1157 game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1 vccd1
+ vccd1 _03770_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13797__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12100__B net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout915_A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_X net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_60_clk_X clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1278_X net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09458_ net1086 _03237_ game.CPU.applesa.ab.absxs.body_x\[68\] net912 vssd1 vssd1
+ vccd1 vccd1 _03701_ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19760__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16735__A2 _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Left_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ net1154 game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1 vccd1
+ vccd1 _03632_ sky130_fd_sc_hd__xor2_1
XANTENNA__12757__A0 _06627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ net798 net315 vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_152_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09622__B1 _03381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_301_Left_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11351_ game.CPU.applesa.ab.check_walls.above.walls\[137\] net769 vssd1 vssd1 vccd1
+ vccd1 _05240_ sky130_fd_sc_hd__xor2_1
XFILLER_0_144_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16523__A _02280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11980__A1 game.CPU.applesa.ab.check_walls.above.walls\[151\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ _04482_ _04484_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__and2_1
X_14070_ net961 game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 _07944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11282_ _05108_ _05113_ _05114_ _05149_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__or4b_1
XFILLER_0_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13358__S net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ net506 _06865_ _06866_ _06572_ net685 vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__o221a_1
XANTENNA__11667__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09925__A1 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13721__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ game.CPU.applesa.ab.count_luck\[4\] game.CPU.applesa.ab.count_luck\[3\] _04420_
+ _04424_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__a31o_1
XANTENNA__15139__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12115__X _06002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14043__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10535__A2 _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__B2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1002 net1003 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__buf_2
XFILLER_0_100_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10164_ _03527_ _04338_ _04340_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__or3_1
Xfanout1013 net1019 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__buf_2
XANTENNA__16120__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1024 net1025 vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_4
XANTENNA__18708__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1035 net1037 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13882__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16671__B2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15426__X _01454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17354__A _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1046 net1051 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_273_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1057 net1058 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__buf_2
X_14972_ net1225 net1252 game.CPU.applesa.ab.check_walls.above.walls\[0\] vssd1 vssd1
+ vccd1 vccd1 _00276_ sky130_fd_sc_hd__and3_1
X_10095_ game.CPU.applesa.twoapples.count_luck\[5\] game.CPU.applesa.twoapples.count_luck\[4\]
+ _04302_ game.CPU.applesa.twoapples.count_luck\[6\] game.CPU.applesa.twoapples.count_luck\[7\]
+ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__a311o_1
X_17760_ game.CPU.applesa.twoapples.count_luck\[3\] game.CPU.applesa.twoapples.count_luck\[2\]
+ _03113_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_163_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1068 game.CPU.applesa.x\[1\] vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_13_clk_X clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1079 game.CPU.bad_collision vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_4
X_16711_ game.writer.tracker.frame\[151\] _02570_ vssd1 vssd1 vccd1 vccd1 _02571_
+ sky130_fd_sc_hd__and2_1
X_13923_ net877 game.CPU.applesa.ab.check_walls.above.walls\[154\] game.CPU.applesa.ab.check_walls.above.walls\[158\]
+ net852 _07792_ vssd1 vssd1 vccd1 vccd1 _07797_ sky130_fd_sc_hd__a221o_1
XANTENNA__17215__A3 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17691_ net1931 _03071_ _03062_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_233_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19290__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19430_ clknet_leaf_41_clk game.writer.tracker.next_frame\[25\] net1352 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[25\] sky130_fd_sc_hd__dfrtp_1
X_16642_ net203 net238 net237 _02290_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__or4_4
XANTENNA__17620__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13854_ game.writer.tracker.frame\[573\] net835 net286 _07724_ vssd1 vssd1 vccd1
+ vccd1 _07728_ sky130_fd_sc_hd__o211a_1
XANTENNA__19966__RESET_B net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18858__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16974__A2 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14434__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ game.writer.tracker.frame\[332\] game.writer.tracker.frame\[333\] net999
+ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16573_ net1757 _02495_ _02496_ net127 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[87\]
+ sky130_fd_sc_hd__a22o_1
X_19361_ clknet_leaf_68_clk _01367_ _00942_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_347_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13785_ net231 _07653_ _07658_ net280 vssd1 vssd1 vccd1 vccd1 _07659_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_28_clk_X clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10997_ _03310_ net404 vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_328_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15524_ _07918_ _01545_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_44_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18312_ net620 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
X_12736_ _06607_ _06608_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__xor2_4
X_19292_ clknet_leaf_71_clk _01336_ _00911_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.steady\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16726__A2 _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18243_ net649 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
X_15455_ _01481_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ _06455_ _06487_ _06493_ _06543_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.absxs.collision
+ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_174_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12748__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14406_ game.CPU.applesa.ab.absxs.body_y\[47\] net942 vssd1 vssd1 vccd1 vccd1 _08280_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_203_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11618_ game.CPU.applesa.ab.check_walls.above.walls\[186\] net765 vssd1 vssd1 vccd1
+ vccd1 _05507_ sky130_fd_sc_hd__xor2_2
X_18174_ net603 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_116_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15386_ _08903_ _08913_ vssd1 vssd1 vccd1 vccd1 _08928_ sky130_fd_sc_hd__or2_1
XANTENNA__15040__C game.CPU.applesa.ab.check_walls.above.walls\[68\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12598_ _06338_ _06339_ _06473_ _06474_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__or4_1
XFILLER_0_142_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17125_ _02379_ net76 net557 vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14337_ _03243_ net1046 net860 game.CPU.applesa.ab.absxs.body_y\[39\] vssd1 vssd1
+ vccd1 vccd1 _08211_ sky130_fd_sc_hd__o22a_1
X_11549_ game.CPU.applesa.ab.check_walls.above.walls\[149\] net314 net258 net789 vssd1
+ vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__16433__A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold507 game.CPU.clock1.counter\[5\] vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold518 game.writer.tracker.frame\[341\] vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10774__A2 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17056_ _02424_ net84 _02687_ net1761 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[379\]
+ sky130_fd_sc_hd__a22o_1
Xhold529 game.CPU.kyle.L1.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14268_ game.CPU.applesa.ab.absxs.body_x\[51\] net874 net962 _03341_ vssd1 vssd1
+ vccd1 vccd1 _08142_ sky130_fd_sc_hd__a22o_1
XANTENNA__13173__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16007_ _02015_ _02016_ _02017_ _02018_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13219_ _07091_ _07092_ net495 vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__mux2_1
XANTENNA__15049__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11988__A2_N net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199_ game.CPU.applesa.ab.absxs.body_x\[66\] net1058 vssd1 vssd1 vccd1 vccd1 _08073_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_55_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_263_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11723__B2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_295_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16111__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15991__B net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16662__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19633__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_185_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12900__S net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17958_ net647 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_302_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09334__X _03577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16909_ _02484_ net95 _02645_ net1669 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[274\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14166__A_N _08028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19252__Q game.CPU.randy.counter1.count\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14400__B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17889_ net614 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__inv_2
XFILLER_0_205_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19628_ clknet_leaf_27_clk game.writer.tracker.next_frame\[223\] net1316 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[223\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13228__A1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19783__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19559_ clknet_leaf_36_clk game.writer.tracker.next_frame\[154\] net1351 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[154\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_200_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16167__X _02179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16608__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_274_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09312_ net1112 game.CPU.applesa.ab.absxs.body_x\[64\] vssd1 vssd1 vccd1 vccd1 _03555_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__16717__A2 _02341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_216_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16327__B net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09510__A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_196_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09243_ game.CPU.applesa.out_random_2\[2\] vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__inv_2
XANTENNA__10462__A1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout231_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12739__B1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09174_ game.CPU.applesa.ab.check_walls.above.walls\[80\] vssd1 vssd1 vccd1 vccd1
+ _03423_ sky130_fd_sc_hd__inv_2
XANTENNA__12834__S0 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16614__Y _02524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13951__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1140_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17142__A2 _02693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout117_X net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19163__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__A2 _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1238_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11962__B2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17158__B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16062__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout698_A net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput16 net16 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_339_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_285_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput38 net38 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_227_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout865_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16653__B2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13467__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14150__X _08024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ game.CPU.apple_location\[6\] vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__inv_2
XANTENNA__11934__B net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16405__B2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17902__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ net546 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.next_head\[3\] sky130_fd_sc_hd__inv_2
XANTENNA__12111__A game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16956__A2 _02413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_316_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10851_ _04748_ _04753_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_296_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout918_X net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13570_ _07442_ _07443_ net501 vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_238_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10782_ game.CPU.applesa.ab.absxs.body_y\[57\] net327 _04722_ net933 vssd1 vssd1
+ vccd1 vccd1 _01008_ sky130_fd_sc_hd__a22o_1
XANTENNA__12442__A2 game.CPU.applesa.twoapples.absxs.next_head\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12521_ game.CPU.applesa.ab.absxs.body_x\[70\] net372 vssd1 vssd1 vccd1 vccd1 _06398_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__15141__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14038__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15240_ game.CPU.kyle.L1.cnt_500hz\[0\] game.CPU.kyle.L1.cnt_500hz\[1\] game.CPU.kyle.L1.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _08801_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19506__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14195__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12452_ game.CPU.applesa.ab.absxs.body_y\[50\] net519 vssd1 vssd1 vccd1 vccd1 _06329_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_191_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11403_ net807 net253 _05291_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_352_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15171_ net1226 net1253 game.CPU.walls.rand_wall.y_final\[3\] vssd1 vssd1 vccd1 vccd1
+ _00265_ sky130_fd_sc_hd__and3_1
X_12383_ game.CPU.applesa.ab.absxs.body_y\[17\] net526 vssd1 vssd1 vccd1 vccd1 _06260_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__17133__A2 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14122_ net879 game.CPU.applesa.ab.check_walls.above.walls\[26\] _03394_ net965 vssd1
+ vssd1 vccd1 vccd1 _07996_ sky130_fd_sc_hd__o22a_1
XFILLER_0_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_327_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11334_ game.CPU.applesa.ab.check_walls.above.walls\[83\] net762 vssd1 vssd1 vccd1
+ vccd1 _05223_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17068__B net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19656__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_249_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16892__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ net1062 _03484_ _03487_ net939 _07920_ vssd1 vssd1 vccd1 vccd1 _07927_ sky130_fd_sc_hd__a221o_1
X_18930_ clknet_leaf_5_clk net1389 _00614_ vssd1 vssd1 vccd1 vccd1 game.CPU.start_pause_button1.eD1.Q1
+ sky130_fd_sc_hd__dfrtp_1
X_11265_ game.CPU.applesa.ab.absxs.body_x\[100\] net415 net402 _03293_ vssd1 vssd1
+ vccd1 vccd1 _05155_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_249_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10508__A2 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11705__A1 game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ game.writer.tracker.frame\[564\] game.writer.tracker.frame\[565\] net1021
+ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__mux2_1
X_10216_ _04386_ _04387_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__xor2_1
X_18861_ clknet_leaf_1_clk _01252_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11196_ _03317_ net534 vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_281_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_280_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_265_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17812_ net182 vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__inv_2
X_10147_ game.CPU.randy.f1.c1.max_i\[1\] _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__or2_1
XFILLER_0_261_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18792_ clknet_leaf_8_clk _01207_ _00529_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[4\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__18680__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17743_ _03102_ _03103_ _03105_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__and3_1
X_14955_ game.CPU.walls.rand_wall.count_luck\[2\] game.CPU.walls.rand_wall.count_luck\[0\]
+ _08730_ game.CPU.walls.rand_wall.count_luck\[1\] vssd1 vssd1 vccd1 vccd1 _08732_
+ sky130_fd_sc_hd__or4b_1
XANTENNA__11844__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10078_ _04213_ _04285_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_50_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13906_ net1069 game.CPU.applesa.ab.check_walls.above.walls\[120\] vssd1 vssd1 vccd1
+ vccd1 _07780_ sky130_fd_sc_hd__or2_1
X_17674_ _03060_ _03061_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__and2b_2
X_14886_ net1125 _08430_ vssd1 vssd1 vccd1 vccd1 _08663_ sky130_fd_sc_hd__and2_1
XANTENNA__15035__C net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_338_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16947__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19413_ clknet_leaf_48_clk game.writer.tracker.next_frame\[8\] net1295 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[8\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19036__CLK net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13837_ game.writer.tracker.frame\[513\] game.writer.tracker.frame\[515\] game.writer.tracker.frame\[516\]
+ game.writer.tracker.frame\[514\] net971 net1008 vssd1 vssd1 vccd1 vccd1 _07711_
+ sky130_fd_sc_hd__mux4_1
X_16625_ net184 _02530_ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__or2_1
XFILLER_0_186_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_348_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_207_Left_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_351_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16556_ _02403_ net144 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__nor2_2
X_19344_ clknet_leaf_72_clk _01359_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.count\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_13768_ game.writer.tracker.frame\[186\] net844 net839 game.writer.tracker.frame\[185\]
+ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__o22a_1
XANTENNA__12433__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16147__B net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ net990 net865 vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__nor2_2
X_15507_ _08404_ _01471_ _01525_ _01529_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__o211a_1
XANTENNA__15051__B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16487_ net168 _02434_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__and2_4
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_19275_ clknet_leaf_7_clk _00045_ _00905_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_13699_ net226 _07572_ _07569_ net284 vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__o211a_1
XANTENNA__19186__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_216_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15438_ _08879_ _08933_ net576 _01465_ vssd1 vssd1 vccd1 vccd1 game.dcx sky130_fd_sc_hd__a22o_1
X_18226_ net664 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14186__A2 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15986__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_300_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15369_ _08905_ _08910_ vssd1 vssd1 vccd1 vccd1 _08911_ sky130_fd_sc_hd__and2b_1
XFILLER_0_142_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18157_ net635 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__inv_2
XANTENNA__13933__A2 game.CPU.applesa.ab.check_walls.above.walls\[35\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17124__A2 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_269_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10747__A2 game.CPU.applesa.ab.absxs.body_y\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_349_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17108_ net161 _02351_ net81 net559 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a31oi_2
Xhold304 game.writer.tracker.frame\[232\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_211_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold315 game.writer.tracker.frame\[264\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
X_18088_ net634 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__inv_2
XFILLER_0_312_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold326 game.writer.tracker.frame\[484\] vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_216_Left_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold337 game.writer.tracker.frame\[573\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 game.writer.tracker.frame\[477\] vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
X_17039_ net188 _02391_ net88 _02683_ net1591 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[366\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_133_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09930_ net1109 net1262 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold359 game.writer.tracker.frame\[179\] vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20050_ game.CPU.en vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
Xfanout806 game.CPU.applesa.ab.check_walls.above.walls\[93\] vssd1 vssd1 vccd1 vccd1
+ net806 sky130_fd_sc_hd__clkbuf_4
X_09861_ net1140 _03309_ _03311_ net1160 _04101_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__a221o_1
Xfanout817 game.CPU.applesa.ab.check_walls.above.walls\[60\] vssd1 vssd1 vccd1 vccd1
+ net817 sky130_fd_sc_hd__buf_2
Xfanout828 game.CPU.applesa.ab.check_walls.above.walls\[22\] vssd1 vssd1 vccd1 vccd1
+ net828 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_284_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout839 net840 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_237_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload16_A clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13449__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09792_ net1133 game.CPU.applesa.ab.absxs.body_y\[43\] vssd1 vssd1 vccd1 vccd1 _04035_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout279_A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16399__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_222_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_225_Left_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_198_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16938__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17060__A1 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10683__A1 game.CPU.applesa.ab.absxs.body_x\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19710__Q game.writer.tracker.frame\[305\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1090_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16338__A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13314__X _07188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19529__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12585__B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_319_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_307_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10386__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout613_A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout234_X net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09226_ game.CPU.applesa.ab.check_walls.above.walls\[176\] vssd1 vssd1 vccd1 vccd1
+ _03475_ sky130_fd_sc_hd__inv_2
XANTENNA__14177__A2 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16571__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15896__B net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19679__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18553__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09157_ game.CPU.applesa.ab.check_walls.above.walls\[49\] vssd1 vssd1 vccd1 vccd1
+ _03406_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_234_Left_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_233_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1143_X net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10738__A2 _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09088_ game.CPU.applesa.ab.absxs.body_y\[59\] vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14305__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16874__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12106__A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout94_A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11050_ _03254_ net322 vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_247_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout868_X net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__A2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16626__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10001_ game.CPU.applesa.twoapples.start_enable game.CPU.applesa.good_collision2
+ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__or2_1
XANTENNA__10271__D game.CPU.applesa.ab.apple_possible\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_322_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15661__A1_N net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11664__B net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09415__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15136__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19059__CLK net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14740_ game.CPU.randy.counter1.count1\[12\] _08565_ vssd1 vssd1 vccd1 vccd1 _08568_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_235_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11952_ net569 _05301_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16929__A2 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17051__A1 _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16519__Y _02460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17051__B2 game.writer.tracker.frame\[375\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10903_ game.CPU.applesa.ab.check_walls.collision_left game.CPU.applesa.ab.check_walls.collision_right
+ _04802_ _04804_ _04791_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__o32a_1
X_14671_ game.CPU.randy.counter1.count1\[5\] _08501_ _08508_ _08509_ vssd1 vssd1 vccd1
+ vccd1 _08510_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_86_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ net828 net302 vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__nand2_1
XANTENNA__16248__A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16410_ _02301_ _02372_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__nor2_4
XANTENNA__13371__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13622_ game.writer.tracker.frame\[273\] game.writer.tracker.frame\[275\] game.writer.tracker.frame\[276\]
+ game.writer.tracker.frame\[274\] net975 net1025 vssd1 vssd1 vccd1 vccd1 _07496_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__15152__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10834_ game.CPU.speed1.Qa\[2\] net1275 _04736_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__mux2_1
X_17390_ _02772_ _02817_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12495__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16341_ net2016 net734 _02329_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[22\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__09150__A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13553_ game.writer.tracker.frame\[69\] game.writer.tracker.frame\[71\] game.writer.tracker.frame\[72\]
+ game.writer.tracker.frame\[70\] net978 net1026 vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10765_ game.CPU.applesa.ab.absxs.body_y\[83\] _04673_ _04674_ game.CPU.applesa.ab.absxs.body_y\[79\]
+ vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14991__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_333_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_325_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12504_ game.CPU.applesa.ab.absxs.body_x\[63\] net530 vssd1 vssd1 vccd1 vccd1 _06381_
+ sky130_fd_sc_hd__xnor2_1
X_19060_ net1191 _00094_ _00731_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[105\]
+ sky130_fd_sc_hd__dfrtp_4
X_16272_ _02274_ net130 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__nand2_4
X_13484_ _07048_ _07131_ _07133_ _07132_ net508 net700 vssd1 vssd1 vccd1 vccd1 _07358_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_171_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10696_ game.CPU.applesa.ab.absxs.body_y\[86\] _04610_ _04611_ game.CPU.applesa.ab.absxs.body_y\[82\]
+ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15223_ game.CPU.applesa.normal1.number\[5\] _08783_ vssd1 vssd1 vccd1 vccd1 _08788_
+ sky130_fd_sc_hd__or2_1
X_18011_ net648 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__inv_2
XFILLER_0_340_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12435_ _06304_ _06306_ _06309_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__or4_1
XANTENNA__17106__A2 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11926__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11926__B2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16414__C _02382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15154_ net1214 net1239 game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1
+ vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16314__B1 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12366_ _06236_ _06237_ _06238_ _06242_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__or4b_1
XFILLER_0_239_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19067__Q game.CPU.applesa.ab.check_walls.above.walls\[112\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16865__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14105_ net1064 game.CPU.applesa.ab.check_walls.above.walls\[49\] vssd1 vssd1 vccd1
+ vccd1 _07979_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11317_ net563 _05192_ game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1 vccd1
+ vccd1 _05206_ sky130_fd_sc_hd__o21a_2
X_19962_ clknet_leaf_43_clk game.writer.tracker.next_frame\[557\] net1306 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[557\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15085_ net1206 net1232 game.CPU.applesa.ab.check_walls.above.walls\[113\] vssd1
+ vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__and3_1
XANTENNA__16270__X _02276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12297_ net828 net420 vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__xnor2_1
X_14036_ net881 game.CPU.applesa.ab.check_walls.above.walls\[113\] game.CPU.applesa.ab.check_walls.above.walls\[115\]
+ net876 vssd1 vssd1 vccd1 vccd1 _07910_ sky130_fd_sc_hd__a22o_1
X_18913_ clknet_leaf_3_clk _00011_ _00597_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.enable_in2
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_52_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11248_ _03226_ net324 vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_276_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19893_ clknet_leaf_28_clk game.writer.tracker.next_frame\[488\] net1309 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[488\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_169_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16617__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18844_ clknet_leaf_0_clk _01235_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_276_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11179_ _05065_ _05066_ _05067_ _05068_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_281_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_182_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19910__RESET_B net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18775_ clknet_leaf_64_clk _01192_ _00512_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[85\]
+ sky130_fd_sc_hd__dfrtp_4
X_15987_ game.CPU.applesa.ab.check_walls.above.walls\[69\] net337 vssd1 vssd1 vccd1
+ vccd1 _01999_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13300__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17726_ _03085_ _03093_ _03094_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__nor3_1
XFILLER_0_166_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14938_ _08664_ _08683_ _08706_ vssd1 vssd1 vccd1 vccd1 _08715_ sky130_fd_sc_hd__or3_1
XFILLER_0_54_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16429__Y _02393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17042__A1 _02535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17657_ net194 _03049_ _03050_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__and3_1
X_14869_ game.CPU.randy.f1.c1.count\[16\] _08653_ net1918 vssd1 vssd1 vccd1 vccd1
+ _08656_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_175_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15062__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16608_ net189 net221 vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__nand2_2
XFILLER_0_9_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17588_ _03004_ _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__or2_2
XFILLER_0_92_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_271_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09060__A game.CPU.applesa.ab.absxs.body_y\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_9_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19327_ clknet_leaf_72_clk net1425 _00932_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twomode.number\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18576__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16539_ net1707 _02469_ _02472_ net124 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[77\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19821__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_311_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18373__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14159__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19258_ clknet_leaf_57_clk _01326_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.count_luck\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_135_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_332_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13367__B1 _07239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16605__B _02480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09011_ game.CPU.applesa.ab.absxs.body_x\[99\] vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18209_ net667 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19189_ clknet_leaf_54_clk net271 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.x_final\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10934__A game.CPU.applesa.ab.absxs.body_x\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_289_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11917__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14406__A game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_331_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11917__B2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold101 game.writer.tracker.frame\[362\] vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 game.writer.tracker.frame\[492\] vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 game.writer.tracker.frame\[226\] vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold134 game.writer.tracker.frame\[326\] vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_257_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 game.writer.tracker.frame\[67\] vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_269_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold156 game.writer.tracker.frame\[250\] vssd1 vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold167 game.writer.tracker.frame\[164\] vssd1 vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_282_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold178 game.writer.tracker.frame\[261\] vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _04152_ _04153_ _04154_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__o21ai_1
Xhold189 game.CPU.applesa.ab.count_luck\[0\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 net604 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__buf_2
XANTENNA__14331__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_300_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_257_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout614 net624 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_4
XANTENNA__19201__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout396_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout625 _08799_ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_298_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20033_ net1381 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 net640 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__buf_4
X_09844_ net924 game.CPU.applesa.ab.absxs.body_x\[31\] game.CPU.applesa.ab.absxs.body_y\[29\]
+ net898 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__o22a_1
Xfanout647 net648 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__buf_4
XFILLER_0_244_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout658 net670 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1103_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 net670 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_2
XANTENNA__17281__A1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11484__B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ net897 game.CPU.applesa.ab.YMAX\[1\] net1170 net902 _04017_ vssd1 vssd1 vccd1
+ vccd1 _04018_ sky130_fd_sc_hd__o221a_1
XANTENNA__14095__A1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout563_A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout184_X net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14095__B2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13980__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19351__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17569__C1 _00293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17033__A1 _02533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10656__A1 game.CPU.applesa.ab.absxs.body_x\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout730_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18919__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_X net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_352_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_293_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_238_Right_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_235_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12883__X _06757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16355__X _02340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18283__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10550_ game.CPU.applesa.ab.absxs.body_x\[31\] net330 _04648_ net930 vssd1 vssd1
+ vccd1 vccd1 _01166_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_242_Left_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09209_ net790 vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10481_ _04176_ _04607_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__nor2_2
XANTENNA__11908__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12220_ net831 net424 vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__nor2_1
XFILLER_0_301_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11659__B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10563__B _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout985_X net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14035__B net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12151_ net792 net386 vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16090__X _02102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout97_X net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11102_ _03225_ net321 vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_246_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12082_ _05350_ _05351_ _05353_ _05355_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__nand4b_1
XANTENNA__16250__B _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15910_ game.CPU.applesa.ab.absxs.body_y\[59\] net435 vssd1 vssd1 vccd1 vccd1 _01922_
+ sky130_fd_sc_hd__xnor2_1
X_11033_ game.CPU.applesa.ab.absxs.body_x\[66\] net410 vssd1 vssd1 vccd1 vccd1 _04923_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__15147__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_251_Left_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16890_ _02267_ net93 _02639_ net1563 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[261\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17272__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__A game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__B net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15841_ _03389_ net337 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15822__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12097__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18560_ clknet_leaf_8_clk _00980_ _00297_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_12984_ _06841_ _06857_ _06639_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__a21o_1
X_15772_ game.CPU.applesa.ab.absxs.body_y\[107\] net435 vssd1 vssd1 vccd1 vccd1 _01784_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__16249__Y _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09432__X _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17511_ _02917_ _02939_ _02938_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__a21o_1
X_11935_ game.CPU.applesa.ab.check_walls.above.walls\[165\] net306 vssd1 vssd1 vccd1
+ vccd1 _05823_ sky130_fd_sc_hd__nand2_1
XANTENNA__18599__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14723_ _08555_ _08556_ net54 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_335_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18491_ net588 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__inv_2
XANTENNA__19844__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17442_ net1258 _02772_ _02827_ _02871_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__a31o_1
XANTENNA__14389__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14654_ game.CPU.randy.counter1.count1\[17\] _08492_ vssd1 vssd1 vccd1 vccd1 _08493_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_358_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13046__C1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11866_ net832 net395 _05753_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_318_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16783__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_257_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13597__B1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13605_ net200 _07478_ net276 vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_205_Right_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10817_ net936 game.CPU.applesa.ab.absxs.body_y\[112\] net233 _04732_ vssd1 vssd1
+ vccd1 vccd1 _00983_ sky130_fd_sc_hd__a31o_1
X_14585_ game.CPU.speed1.Qa\[2\] _03520_ _08446_ vssd1 vssd1 vccd1 vccd1 _08447_ sky130_fd_sc_hd__o21ai_1
X_17373_ net1117 _02802_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__or2_1
X_11797_ net749 _05441_ _05440_ net575 vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__18193__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19112_ net1180 _00151_ _00783_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[157\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10457__C _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13536_ game.writer.tracker.frame\[85\] game.writer.tracker.frame\[87\] game.writer.tracker.frame\[88\]
+ game.writer.tracker.frame\[86\] net978 net1028 vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__mux4_1
X_16324_ net196 _02315_ _02317_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__o21a_2
XANTENNA__16535__B1 _02470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ game.CPU.applesa.ab.absxs.body_y\[115\] _04663_ _04664_ game.CPU.applesa.ab.absxs.body_y\[111\]
+ vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19994__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13349__A0 _06627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_314_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16255_ net872 _08028_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__or2_1
X_19043_ net1191 _00274_ _00714_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[88\]
+ sky130_fd_sc_hd__dfrtp_4
X_13467_ net214 _07340_ _07337_ net285 vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__a211o_1
XANTENNA__11252__A1_N game.CPU.applesa.ab.absxs.body_x\[115\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10679_ net936 game.CPU.applesa.ab.absxs.body_x\[112\] net233 _04706_ vssd1 vssd1
+ vccd1 vccd1 _01095_ sky130_fd_sc_hd__a31o_1
XFILLER_0_125_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ game.CPU.applesa.normal1.number\[2\] _08768_ vssd1 vssd1 vccd1 vccd1 _08774_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12021__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12418_ game.CPU.applesa.ab.absxs.body_x\[34\] net374 vssd1 vssd1 vccd1 vccd1 _06295_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09568__A2 game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16186_ game.CPU.applesa.ab.check_walls.above.walls\[105\] net475 net466 game.CPU.applesa.ab.check_walls.above.walls\[106\]
+ _01680_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__a221o_1
X_13398_ _06876_ _06889_ net685 vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_346_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19224__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15137_ net1209 net1234 game.CPU.applesa.ab.check_walls.above.walls\[165\] vssd1
+ vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17537__A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12349_ game.CPU.applesa.ab.absxs.body_x\[39\] net529 net527 game.CPU.applesa.ab.absxs.body_y\[37\]
+ _06225_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_130_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19945_ clknet_leaf_38_clk game.writer.tracker.next_frame\[540\] net1324 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[540\] sky130_fd_sc_hd__dfrtp_1
X_15068_ net1212 net1238 game.CPU.applesa.ab.check_walls.above.walls\[96\] vssd1 vssd1
+ vccd1 vccd1 _00093_ sky130_fd_sc_hd__and3_1
XANTENNA__13276__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13521__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14019_ net1062 _03480_ _03481_ net984 _07890_ vssd1 vssd1 vccd1 vccd1 _07893_ sky130_fd_sc_hd__a221o_1
XANTENNA__15057__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_339_Left_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19876_ clknet_leaf_27_clk game.writer.tracker.next_frame\[471\] net1316 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[471\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_226_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19374__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17263__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10886__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18827_ clknet_leaf_1_clk _01218_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__dfxtp_1
XANTENNA__10886__B2 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14077__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14077__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15813__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ net1087 _03238_ _03239_ net1104 _03802_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__a221o_1
XFILLER_0_207_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18758_ clknet_leaf_12_clk _01175_ _00495_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[52\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_108_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12627__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_357_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17709_ net758 game.CPU.applesa.normal1.counter_normal vssd1 vssd1 vccd1 vccd1 _01320_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_349_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11835__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09491_ net915 game.CPU.applesa.ab.check_walls.above.walls\[185\] game.CPU.applesa.ab.check_walls.above.walls\[189\]
+ net898 _03733_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__a221o_1
X_18689_ clknet_leaf_62_clk _01106_ _00426_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10929__A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_349_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13037__C1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11835__A1_N net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13588__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16175__X _02187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13683__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16616__A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19349__D net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout311_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1053_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_320_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_230_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16829__B2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13760__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13975__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1220_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1318_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19717__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15238__Y _00293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout680_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 _04817_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10670__Y _04701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16070__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout411 _04812_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_4
XFILLER_0_347_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13512__B1 _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 net424 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout778_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout433 net436 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_8
Xfanout444 _08427_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1106_X net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17254__A1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout466 net470 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_4
XANTENNA__16057__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout477 net478 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_4
X_09827_ net1159 game.CPU.applesa.ab.absxs.body_y\[12\] vssd1 vssd1 vccd1 vccd1 _04070_
+ sky130_fd_sc_hd__or2_1
X_20016_ net1277 vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_232_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout488 net489 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_307_Right_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12878__X _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout499 _06596_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout945_A net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18741__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19867__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09758_ net1086 game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1 vccd1
+ vccd1 _04001_ sky130_fd_sc_hd__nand2_1
XANTENNA__12618__A2 game.CPU.applesa.twoapples.absxs.next_head\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_241_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17006__A1 _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout57_A _02692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ net1092 game.CPU.applesa.ab.absxs.body_x\[6\] vssd1 vssd1 vccd1 vccd1 _03932_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_185_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09537__A2_N net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ _05599_ _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__nand2_1
XANTENNA__17910__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13579__B1 _07452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout900_X net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11651_ game.CPU.applesa.ab.check_walls.above.walls\[11\] net764 vssd1 vssd1 vccd1
+ vccd1 _05540_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_154_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16526__A _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14240__B2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16780__A3 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout62 net65 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_2
XANTENNA__14972__C game.CPU.applesa.ab.check_walls.above.walls\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10602_ net1268 _04590_ net329 game.CPU.applesa.ab.absxs.body_x\[87\] vssd1 vssd1
+ vccd1 vccd1 _01138_ sky130_fd_sc_hd__a22o_1
XFILLER_0_308_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14370_ game.CPU.applesa.ab.absxs.body_y\[118\] net953 vssd1 vssd1 vccd1 vccd1 _08244_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__16517__B1 _02458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout73 net74 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_2
X_11582_ _05454_ _05470_ _05457_ _05466_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__or4b_2
Xfanout84 net85 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_330_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout95 net97 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_2
X_13321_ net510 _06709_ net703 vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10533_ net849 _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_21_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10801__B2 game.CPU.applesa.ab.absxs.body_y\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14046__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ game.CPU.applesa.ab.absxs.body_x\[46\] net468 vssd1 vssd1 vccd1 vccd1 _02052_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ _07124_ _07125_ net508 vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__mux2_1
XANTENNA__11389__B net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ net932 game.CPU.applesa.ab.absxs.body_x\[98\] _04594_ _04597_ vssd1 vssd1
+ vccd1 vccd1 _01201_ sky130_fd_sc_hd__a31o_1
X_12203_ game.CPU.applesa.ab.check_walls.above.walls\[198\] net418 vssd1 vssd1 vccd1
+ vccd1 _06089_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_295_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13885__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13183_ _07053_ _07054_ _07056_ _07055_ net497 net689 vssd1 vssd1 vccd1 vccd1 _07057_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__16261__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10395_ _04537_ _04540_ _04546_ game.CPU.applesa.ab.good_collision _03191_ vssd1
+ vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_94_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19397__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ net815 net389 vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_36_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17991_ net640 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__inv_2
XFILLER_0_236_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13096__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19730_ clknet_leaf_19_clk game.writer.tracker.next_frame\[325\] net1342 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[325\] sky130_fd_sc_hd__dfrtp_1
X_16942_ _02299_ net163 net87 _02653_ net1590 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[299\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12065_ game.CPU.applesa.ab.check_walls.above.walls\[127\] net294 net288 net794 vssd1
+ vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_341_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17245__A1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ _04897_ _04900_ _04901_ _04905_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__or4_1
X_19661_ clknet_leaf_23_clk game.writer.tracker.next_frame\[256\] net1344 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[256\] sky130_fd_sc_hd__dfrtp_1
X_16873_ _02551_ net108 _02629_ net1665 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[254\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14059__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14059__B2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18612_ clknet_leaf_63_clk _01029_ _00349_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[98\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_189_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15824_ game.CPU.applesa.ab.absxs.body_y\[91\] net431 net449 game.CPU.applesa.ab.absxs.body_y\[88\]
+ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__o2bb2a_1
X_19592_ clknet_leaf_37_clk game.writer.tracker.next_frame\[187\] net1355 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[187\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12609__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_148_Left_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18543_ net611 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__inv_2
X_12967_ net240 _06827_ _06832_ _06840_ net189 vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__a311o_1
X_15755_ game.CPU.applesa.ab.check_walls.above.walls\[5\] net447 vssd1 vssd1 vccd1
+ vccd1 _01767_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16205__C1 _02210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09486__B2 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ net829 net313 net308 net830 vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__o22ai_1
X_14706_ _04486_ _08544_ vssd1 vssd1 vccd1 vccd1 _08545_ sky130_fd_sc_hd__nor2_1
X_18474_ net638 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
X_12898_ _06768_ _06770_ net685 vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15043__C game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15686_ game.CPU.applesa.ab.absxs.body_x\[4\] net273 vssd1 vssd1 vccd1 vccd1 _01698_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_346_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17425_ net846 net428 _02825_ _02854_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a31o_1
X_14637_ game.CPU.clock1.counter\[18\] _08479_ net267 vssd1 vssd1 vccd1 vccd1 _08481_
+ sky130_fd_sc_hd__o21ai_1
X_11849_ net751 _05365_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_177_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17356_ _04638_ _02784_ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__nand2_1
X_14568_ game.CPU.start_pause_button1.eD1.Q2 game.CPU.start_pause_button1.eD1.Q1 vssd1
+ vssd1 vccd1 vccd1 _08432_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_129_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16307_ net1995 net720 _02304_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[13\]
+ sky130_fd_sc_hd__and3_1
X_13519_ _07368_ _07369_ net217 vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17287_ net111 _02512_ _02752_ game.writer.tracker.frame\[545\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[545\] sky130_fd_sc_hd__a22o_1
X_14499_ game.CPU.apple_location\[5\] net958 vssd1 vssd1 vccd1 vccd1 _08373_ sky130_fd_sc_hd__nand2_1
XANTENNA__10484__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09600__A1_N net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload10 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 clkload10/X sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_157_Left_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18614__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload21 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_12
X_19026_ net1195 _00256_ _00697_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[71\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_302_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16238_ net507 net835 _02226_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a21o_1
Xclkload32 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__15994__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload43 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload54 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12545__A1 game.CPU.applesa.ab.absxs.body_x\[40\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkload65 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__clkinv_16
XFILLER_0_301_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14243__X _08117_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09410__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16169_ _02154_ _02155_ _02179_ _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__and4_1
XANTENNA__09410__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_266_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_347_Left_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08991_ game.CPU.applesa.ab.absxs.body_x\[55\] vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__inv_2
XANTENNA__14298__A1 game.CPU.applesa.ab.absxs.body_y\[52\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10931__B net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18764__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19928_ clknet_leaf_48_clk game.writer.tracker.next_frame\[523\] net1302 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[523\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17236__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_305_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19859_ clknet_leaf_20_clk game.writer.tracker.next_frame\[454\] net1317 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[454\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_214_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_166_Left_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_317_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09612_ net1102 _03287_ game.CPU.applesa.ab.absxs.body_y\[116\] net893 _03848_ vssd1
+ vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__a221o_1
XFILLER_0_183_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09543_ net914 game.CPU.applesa.ab.XMAX\[1\] net1172 net919 vssd1 vssd1 vccd1 vccd1
+ _03786_ sky130_fd_sc_hd__o22a_1
XANTENNA__11808__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13273__A2 _07144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_203_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout359_A net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11284__A1 _04936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15802__X _01814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_356_Left_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_333_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_277_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09474_ net1147 _03478_ game.CPU.applesa.ab.check_walls.above.walls\[182\] net905
+ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__a22o_1
XANTENNA__12481__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_349_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_219_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_290_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16346__A _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1170_A game.CPU.applesa.ab.YMAX\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout526_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15250__A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload4 clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_8
XPHY_EDGE_ROW_175_Left_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16065__B net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17172__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1056_X net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout895_A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13733__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12813__S net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09401__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14153__X _08027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09401__B2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_258_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10180_ net891 _04369_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_292_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14313__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 net1216 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_243_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17905__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09407__B net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1217 net1218 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__clkbuf_2
Xfanout230 net232 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__buf_4
XANTENNA__15128__C game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1228 game.CPU.walls.rand_wall.start_enable vssd1 vssd1 vccd1 vccd1 net1228
+ sky130_fd_sc_hd__clkbuf_2
Xfanout241 net243 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_4
XANTENNA__17227__A1 _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_184_Left_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1239 net1240 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__clkbuf_2
Xfanout252 net253 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_4
Xfanout263 _04667_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
XANTENNA_fanout850_X net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout274 _06610_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_4
Xfanout285 net286 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_227_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout296 net298 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_2
XANTENNA__11953__A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13870_ net1060 _03370_ _03371_ net1052 vssd1 vssd1 vccd1 vccd1 _07744_ sky130_fd_sc_hd__a22o_1
XANTENNA__16986__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ _06690_ _06691_ _06693_ _06692_ net491 net687 vssd1 vssd1 vccd1 vccd1 _06695_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09423__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15144__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11672__B net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_319_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09468__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09468__B2 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11017__X _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_290_Right_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12752_ _06624_ _06625_ net477 vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__mux2_1
X_15540_ net943 net834 _01527_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_243_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16202__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11703_ _05590_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__nand2_1
X_15471_ _01497_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__inv_2
XANTENNA__10483__C1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12683_ _06556_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_254_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ net68 net143 net120 _02733_ net1616 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[487\]
+ sky130_fd_sc_hd__a32o_1
X_14422_ _03259_ net1067 net859 game.CPU.applesa.ab.absxs.body_y\[111\] _08292_ vssd1
+ vssd1 vccd1 vccd1 _08296_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_193_Left_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15160__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12379__A2_N net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ game.CPU.applesa.ab.check_walls.above.walls\[155\] net761 vssd1 vssd1 vccd1
+ vccd1 _05523_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_139_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18190_ net635 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_343_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12775__A1 game.writer.tracker.frame\[129\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17141_ net185 _02412_ net80 _02714_ net1529 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[437\]
+ sky130_fd_sc_hd__a32o_1
X_14353_ game.CPU.applesa.ab.absxs.body_y\[32\] net869 net857 game.CPU.applesa.ab.absxs.body_y\[35\]
+ _08224_ vssd1 vssd1 vccd1 vccd1 _08227_ sky130_fd_sc_hd__o221a_1
XFILLER_0_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11565_ game.CPU.applesa.ab.check_walls.above.walls\[135\] net258 vssd1 vssd1 vccd1
+ vccd1 _05454_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13304_ game.writer.tracker.frame\[0\] game.writer.tracker.frame\[2\] game.writer.tracker.frame\[3\]
+ game.writer.tracker.frame\[1\] net970 net1002 vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_42_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17072_ _02454_ net59 _02694_ net2012 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[388\]
+ sky130_fd_sc_hd__a22o_1
X_10516_ net1122 _04177_ _04578_ _04620_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__o31a_1
XFILLER_0_296_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14284_ _08155_ _08156_ _08157_ _08154_ vssd1 vssd1 vccd1 vccd1 _08158_ sky130_fd_sc_hd__a211o_1
X_11496_ game.CPU.applesa.ab.check_walls.above.walls\[170\] net766 vssd1 vssd1 vccd1
+ vccd1 _05385_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18787__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_311_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13235_ game.writer.tracker.frame\[480\] game.writer.tracker.frame\[481\] net1011
+ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_268_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16023_ _03230_ net350 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__xnor2_1
X_10447_ net1117 net1121 net1124 net1119 vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_343_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10538__B1 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_311_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_268_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13166_ _07032_ _07034_ net684 vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__mux2_1
XANTENNA__11847__B net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10378_ net1153 game.CPU.apple_location2\[4\] vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__nor2_1
XANTENNA__19075__Q game.CPU.applesa.ab.check_walls.above.walls\[120\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14223__B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12117_ _05968_ _05985_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__or3_1
XANTENNA__13488__C1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13097_ net220 _06970_ net276 vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__a21o_1
XANTENNA__12024__A game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17974_ net643 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__inv_2
XANTENNA__15038__C game.CPU.applesa.ab.check_walls.above.walls\[66\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17218__A1 _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19713_ clknet_leaf_35_clk game.writer.tracker.next_frame\[308\] net1340 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[308\] sky130_fd_sc_hd__dfrtp_1
X_16925_ _02430_ _02644_ _02649_ net1678 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[286\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_264_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12048_ _05568_ _05569_ _05570_ _05572_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_284_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12959__A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11502__A2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19644_ clknet_leaf_15_clk game.writer.tracker.next_frame\[239\] net1289 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[239\] sky130_fd_sc_hd__dfrtp_1
X_16856_ _02541_ net104 _02623_ net2052 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[242\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_284_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12678__B net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16441__A2 net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15807_ _03410_ net271 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__xnor2_1
X_19575_ clknet_leaf_50_clk game.writer.tracker.next_frame\[170\] net1279 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[170\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09459__A1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15054__B net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16787_ _02465_ net104 _02596_ game.writer.tracker.frame\[200\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[200\] sky130_fd_sc_hd__a22o_1
XANTENNA__19412__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09459__B2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_179_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10479__A _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16718__X _02574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13999_ net880 game.CPU.applesa.ab.check_walls.above.walls\[74\] game.CPU.applesa.ab.check_walls.above.walls\[78\]
+ net855 _07868_ vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_354_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18526_ net586 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__inv_2
XANTENNA__11266__A1 game.CPU.applesa.ab.absxs.body_x\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15738_ _03470_ net350 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11266__B2 game.CPU.applesa.ab.absxs.body_y\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_303_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18457_ net654 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15669_ net800 net432 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_334_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15070__A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17408_ net741 _02837_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__nor2_1
X_09190_ net801 vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__inv_2
XANTENNA__19562__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13412__C1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18388_ net599 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_334_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17339_ net1116 _04582_ _08749_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__nor3_1
XANTENNA__17154__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16901__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload46_A clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_287_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_259_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19009_ net1194 _00237_ _00680_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10792__A3 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17711__A_N _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10529__B1 _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout107_A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_307_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_302_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09508__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_227_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08974_ game.CPU.applesa.ab.absxs.body_x\[7\] vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1016_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17209__A1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold16 game.CPU.up_button.eD1.Q1 vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_282_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold27 game.CPU.applesa.off_bc.D vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 game.CPU.applesa.normal1.number\[4\] vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold49 game.CPU.walls.rand_wall.count\[3\] vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13464__S net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_279_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout476_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16968__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16432__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11492__B net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout643_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09526_ net1126 game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1 vccd1
+ vccd1 _03769_ sky130_fd_sc_hd__xor2_1
XANTENNA__17460__A _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12454__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15899__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19905__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09457_ net912 game.CPU.applesa.ab.absxs.body_x\[68\] game.CPU.applesa.ab.absxs.body_y\[68\]
+ net893 vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09870__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09870__B2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_X net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout908_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09388_ net1082 _03467_ game.CPU.applesa.ab.check_walls.above.walls\[165\] net897
+ _03630_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09622__A1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18291__A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09622__B2 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_352_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ net742 _05235_ _05238_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__a21o_1
XFILLER_0_163_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13639__S net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout898_X net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10301_ game.CPU.clock1.game_state\[0\] net1264 vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_61_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11948__A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ game.CPU.applesa.ab.absxs.body_x\[39\] net545 net542 game.CPU.applesa.ab.absxs.body_y\[37\]
+ _05170_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14324__A game.CPU.applesa.ab.absxs.body_x\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_293_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13020_ net697 _06893_ _06892_ vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10232_ game.CPU.applesa.ab.count_luck\[4\] game.CPU.applesa.ab.count_luck\[3\] vssd1
+ vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__nand2_1
XANTENNA__09418__A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15139__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14043__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1003 net1004 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__buf_2
X_10163_ net1078 _03527_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__or2_4
Xfanout1014 net1016 vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__clkbuf_4
Xfanout1025 net1041 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__buf_2
XFILLER_0_218_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1036 net1037 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_4
Xfanout1047 net1051 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_2
X_14971_ _04256_ _08746_ _08747_ _03522_ net1243 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__o32a_1
X_10094_ game.CPU.applesa.twoapples.count_luck\[3\] _04261_ vssd1 vssd1 vccd1 vccd1
+ _04302_ sky130_fd_sc_hd__or2_1
XANTENNA__19435__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1058 net1059 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_163_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1069 net1071 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_4
XANTENNA__13227__X _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16710_ _02491_ net63 _02570_ net1536 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[150\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15155__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13922_ net948 _03462_ net788 net856 _07795_ vssd1 vssd1 vccd1 vccd1 _07796_ sky130_fd_sc_hd__a221o_1
X_17690_ _03062_ _03071_ _03072_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__nor3_1
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12498__B net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16641_ game.writer.tracker.frame\[113\] _02537_ _02538_ net124 vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[113\] sky130_fd_sc_hd__a22o_1
X_13853_ net286 _07721_ _07725_ _07726_ vssd1 vssd1 vccd1 vccd1 _07727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15631__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12804_ game.writer.tracker.frame\[336\] game.writer.tracker.frame\[337\] net1017
+ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__mux2_2
X_19360_ clknet_leaf_69_clk _01366_ _00941_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_16572_ net171 net151 net69 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__and3_2
XANTENNA__19585__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13784_ net216 _07657_ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10996_ game.CPU.applesa.ab.absxs.body_y\[44\] net535 vssd1 vssd1 vccd1 vccd1 _04886_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_347_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09310__B1 game.CPU.applesa.ab.absxs.body_y\[52\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18311_ net621 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
X_15523_ net965 net943 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12735_ _06607_ _06608_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_44_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19291_ clknet_leaf_6_clk _01335_ _00910_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.max_i\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09861__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09861__B2 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18242_ net650 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
XFILLER_0_270_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15454_ _01449_ _01454_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_182_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _06302_ _06392_ _06500_ _06542_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__and4_1
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10746__B net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14405_ _08273_ _08276_ _08277_ _08278_ vssd1 vssd1 vccd1 vccd1 _08279_ sky130_fd_sc_hd__or4_1
X_11617_ game.CPU.applesa.ab.check_walls.above.walls\[189\] net315 vssd1 vssd1 vccd1
+ vccd1 _05506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18173_ net602 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__inv_2
XANTENNA__17136__B1 _02713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15385_ _08899_ _08916_ vssd1 vssd1 vccd1 vccd1 _08927_ sky130_fd_sc_hd__or2_1
X_12597_ game.CPU.applesa.ab.absxs.body_y\[111\] net366 vssd1 vssd1 vccd1 vccd1 _06474_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_116_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17124_ _02378_ net76 _02709_ game.writer.tracker.frame\[425\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[425\] sky130_fd_sc_hd__a22o_1
X_11548_ net789 net258 net314 game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1
+ vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__a2bb2o_1
X_14336_ _08197_ _08198_ _08202_ _08203_ _08209_ vssd1 vssd1 vccd1 vccd1 _08210_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15698__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 game.writer.tracker.frame\[524\] vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11858__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17055_ _02423_ net83 _02687_ net1679 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[378\]
+ sky130_fd_sc_hd__a22o_1
Xhold519 game.writer.tracker.frame\[134\] vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14267_ _08135_ _08140_ vssd1 vssd1 vccd1 vccd1 _08141_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11479_ net777 _05367_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__xor2_1
XANTENNA__14234__A game.CPU.applesa.ab.absxs.body_x\[115\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13173__A1 _06984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13218_ game.writer.tracker.frame\[418\] game.writer.tracker.frame\[419\] net1024
+ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_256_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16006_ game.CPU.applesa.ab.absxs.body_x\[60\] net271 vssd1 vssd1 vccd1 vccd1 _02018_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_0_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15049__B net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14198_ _08069_ _08070_ _08071_ vssd1 vssd1 vccd1 vccd1 _08072_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_55_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12920__A1 _06783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_263_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ game.writer.tracker.frame\[180\] game.writer.tracker.frame\[181\] net1036
+ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16662__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17957_ net647 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
XFILLER_0_252_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_302_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16908_ _02482_ net95 _02645_ game.writer.tracker.frame\[273\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[273\] sky130_fd_sc_hd__a22o_1
X_17888_ net634 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__inv_2
XANTENNA__19928__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19627_ clknet_leaf_26_clk game.writer.tracker.next_frame\[222\] net1316 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[222\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_205_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16839_ _02531_ net98 net715 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__o21a_1
XFILLER_0_164_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13228__A2 _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12201__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19558_ clknet_leaf_36_clk game.writer.tracker.next_frame\[153\] net1349 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[153\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_289_Left_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_200_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09311_ _03547_ _03548_ _03549_ _03551_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__or4_1
X_18509_ net579 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_274_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19489_ clknet_leaf_23_clk game.writer.tracker.next_frame\[84\] net1339 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[84\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18952__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16717__A3 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_216_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09242_ net1404 vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_196_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09173_ game.CPU.applesa.ab.check_walls.above.walls\[76\] vssd1 vssd1 vccd1 vccd1
+ _03422_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_313_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16183__X _02195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16624__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout224_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12834__S1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19357__D game.CPU.applesa.twoapples.absxs.next_head\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18612__Q game.CPU.applesa.ab.absxs.body_y\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_298_Left_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_330_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput17 net17 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_77_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XANTENNA__14361__B1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_285_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput39 net39 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XANTENNA__19458__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_227_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13983__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1300_A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_X net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08957_ game.CPU.apple_location2\[0\] vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout760_A net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13467__A2 _07340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout479_X net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12111__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_224_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16956__A3 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_316_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__inv_2
XFILLER_0_357_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_296_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12978__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_345_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09509_ net1142 game.CPU.applesa.ab.absxs.body_y\[50\] vssd1 vssd1 vccd1 vccd1 _03752_
+ sky130_fd_sc_hd__nand2_1
X_10781_ _03307_ net327 vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_238_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09843__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09843__B2 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12520_ game.CPU.applesa.ab.absxs.body_x\[68\] net383 vssd1 vssd1 vccd1 vccd1 _06397_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11650__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_251_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12451_ game.CPU.applesa.ab.absxs.body_x\[50\] net371 vssd1 vssd1 vccd1 vccd1 _06328_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_352_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11590__A1_N net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16534__A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11402_ net807 net252 _05286_ _05287_ _05290_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_325_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15170_ net1227 net1254 game.CPU.walls.rand_wall.y_final\[2\] vssd1 vssd1 vccd1 vccd1
+ _00254_ sky130_fd_sc_hd__and3_1
XANTENNA__11402__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12382_ game.CPU.applesa.ab.absxs.body_y\[19\] net367 vssd1 vssd1 vccd1 vccd1 _06259_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17133__A3 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13369__S net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14121_ net870 net826 game.CPU.applesa.ab.check_walls.above.walls\[29\] net865 vssd1
+ vssd1 vccd1 vccd1 _07995_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_340_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11333_ _05218_ _05219_ _05220_ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11678__A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_327_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14054__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14052_ net882 game.CPU.applesa.ab.check_walls.above.walls\[193\] _03486_ net984
+ _07925_ vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__a221o_1
XANTENNA__09148__A game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16892__A2 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11397__B net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11264_ game.CPU.applesa.ab.absxs.body_y\[102\] net539 net534 _03295_ _05153_ vssd1
+ vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_249_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14989__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ game.writer.tracker.frame\[568\] game.writer.tracker.frame\[569\] net1021
+ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__mux2_1
XANTENNA__11705__A2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ _04406_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__xnor2_1
X_18860_ clknet_leaf_1_clk _01251_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11195_ game.CPU.applesa.ab.absxs.body_y\[23\] net397 vssd1 vssd1 vccd1 vccd1 _05085_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__08987__A game.CPU.applesa.ab.absxs.body_x\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18825__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17811_ _08934_ _01438_ _03143_ _03145_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__a31o_1
XFILLER_0_206_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10146_ _04338_ _04340_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__nor2_2
XFILLER_0_265_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18791_ clknet_leaf_4_clk _01206_ _00528_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_273_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14501__B net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17742_ game.CPU.applesa.ab.count\[1\] game.CPU.applesa.ab.count\[0\] net1167 game.CPU.applesa.ab.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__a31o_1
XANTENNA__11469__A1 game.CPU.applesa.ab.check_walls.above.walls\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ net910 _04211_ _04212_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__or3b_1
X_14954_ game.CPU.walls.rand_wall.count_luck\[4\] game.CPU.walls.rand_wall.count_luck\[3\]
+ _08725_ _08729_ vssd1 vssd1 vccd1 vccd1 _08731_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_50_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13905_ net1069 game.CPU.applesa.ab.check_walls.above.walls\[120\] vssd1 vssd1 vccd1
+ vccd1 _07779_ sky130_fd_sc_hd__nand2_1
X_17673_ _03362_ _08741_ _08745_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__a21o_1
X_14885_ _08660_ _08661_ vssd1 vssd1 vccd1 vccd1 _08662_ sky130_fd_sc_hd__and2b_1
XANTENNA__18975__CLK net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15604__B1 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_338_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19412_ clknet_leaf_48_clk game.writer.tracker.next_frame\[7\] net1295 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload2_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16624_ net201 _02529_ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__or2_1
X_13836_ net287 _07708_ _07709_ net245 vssd1 vssd1 vccd1 vccd1 _07710_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19343_ clknet_leaf_72_clk _01358_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.count\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16555_ net170 _02403_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__nor2_2
XFILLER_0_97_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13767_ game.writer.tracker.frame\[187\] net711 net675 game.writer.tracker.frame\[188\]
+ vssd1 vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__o22a_1
X_10979_ _03333_ net534 vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__xnor2_1
X_15506_ _01506_ _01524_ _01528_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__or3_1
X_12718_ _06578_ _06590_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__xor2_1
XANTENNA__11641__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19274_ clknet_leaf_7_clk _00044_ _00904_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[14\]
+ sky130_fd_sc_hd__dfrtp_2
X_16486_ net197 _02392_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__nor2_4
X_13698_ _07570_ _07571_ net490 vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__mux2_1
X_18225_ net649 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__inv_2
X_15437_ _01435_ _01457_ _01464_ _01455_ _01461_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12649_ _06275_ _06277_ _06278_ _06279_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__or4_1
XFILLER_0_209_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18156_ net635 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__inv_2
X_15368_ game.writer.updater.commands.cmd_num\[1\] game.writer.updater.commands.cmd_num\[0\]
+ game.writer.updater.commands.cmd_num\[2\] game.writer.updater.commands.cmd_num\[3\]
+ vssd1 vssd1 vccd1 vccd1 _08910_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_130_Left_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17107_ net160 _02348_ net81 _02704_ net1580 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[413\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__13279__S net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10747__A3 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11588__A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_349_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold305 game.writer.tracker.frame\[75\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
X_14319_ game.CPU.applesa.ab.absxs.body_y\[57\] net866 _08188_ _08189_ _08192_ vssd1
+ vssd1 vccd1 vccd1 _08193_ sky130_fd_sc_hd__a221o_1
XANTENNA__19600__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold316 game.writer.tracker.frame\[541\] vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
X_18087_ net634 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__inv_2
X_15299_ net757 _08844_ _08845_ _08846_ _08847_ vssd1 vssd1 vccd1 vccd1 _08848_ sky130_fd_sc_hd__a32o_1
XFILLER_0_123_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold327 game.writer.tracker.frame\[218\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_312_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold338 game.writer.tracker.frame\[78\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold349 game.writer.tracker.frame\[313\] vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
X_17038_ _02238_ _02517_ _02619_ net713 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__o31a_1
XANTENNA__14343__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_309_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_320_Left_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11100__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ _04100_ _04102_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__nand2_1
Xfanout807 game.CPU.applesa.ab.check_walls.above.walls\[92\] vssd1 vssd1 vccd1 vccd1
+ net807 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout818 game.CPU.applesa.ab.check_walls.above.walls\[55\] vssd1 vssd1 vccd1 vccd1
+ net818 sky130_fd_sc_hd__clkbuf_4
Xfanout829 game.CPU.applesa.ab.check_walls.above.walls\[15\] vssd1 vssd1 vccd1 vccd1
+ net829 sky130_fd_sc_hd__clkbuf_4
XANTENNA__19750__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09791_ net1110 game.CPU.applesa.ab.absxs.body_x\[40\] vssd1 vssd1 vccd1 vccd1 _04034_
+ sky130_fd_sc_hd__xnor2_1
X_18989_ net1197 _00215_ _00660_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[34\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10380__A1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10380__B2 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12657__B1 game.CPU.applesa.twoapples.absxs.next_head\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12212__A game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_219_Right_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16399__A1 _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_222_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout174_A _06702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16178__X _02190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13742__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_198_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15523__A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11880__A1 game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09521__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11770__B net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09878__D _04075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A _08429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19130__CLK net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_341_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09225_ game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1 vssd1 vccd1 vccd1
+ _03474_ sky130_fd_sc_hd__inv_2
XANTENNA__13909__B1 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_350_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16571__A1 _02243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16354__A _08028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1250_A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout227_X net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1348_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09589__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_12_clk_X clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ net820 vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_233_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16073__B net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14145__Y _08019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19280__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09087_ game.CPU.applesa.ab.absxs.body_y\[64\] vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1136_X net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14334__B1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16874__A2 _02432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout975_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12106__B net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_X clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11010__B net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11699__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout87_A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10000_ net1162 _03492_ game.CPU.applesa.good_collision2 _03212_ vssd1 vssd1 vccd1
+ vccd1 _01364_ sky130_fd_sc_hd__a211o_1
XANTENNA__16087__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__B net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ game.CPU.apple_location2\[2\] _04208_ _04209_ net1900 vssd1 vssd1 vccd1 vccd1
+ _01375_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_322_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18998__CLK net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17913__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12648__B1 game.CPU.applesa.twoapples.absxs.next_head\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09415__B game.CPU.applesa.ab.absxs.body_y\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13845__C1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15136__C game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _05831_ _05832_ _05835_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout930_X net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13860__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14975__C game.CPU.applesa.ab.check_walls.above.walls\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17051__A2 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10902_ _04778_ _04790_ _04796_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a21oi_1
X_11882_ _05754_ _05758_ _05760_ _05769_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__a31o_1
X_14670_ game.CPU.randy.counter1.count1\[7\] _08498_ vssd1 vssd1 vccd1 vccd1 _08509_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__13299__S1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16248__B net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__A0 _06943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13621_ _07491_ _07494_ net213 vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__mux2_1
X_10833_ net720 vssd1 vssd1 vccd1 vccd1 game.CPU.button_reset_in sky130_fd_sc_hd__inv_2
XANTENNA__15152__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__B net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14049__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09816__A1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09816__B2 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16340_ net2011 net734 _02329_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[21\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_251_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13552_ _07424_ _07425_ net476 vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__mux2_1
X_10764_ game.CPU.applesa.ab.absxs.body_y\[88\] _04590_ net329 game.CPU.applesa.ab.absxs.body_y\[84\]
+ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_333_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12503_ game.CPU.applesa.ab.absxs.body_x\[62\] net373 vssd1 vssd1 vccd1 vccd1 _06380_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13888__A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16271_ _02273_ _02275_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__nor2_1
X_13483_ net226 _07356_ _07353_ net277 vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__a211o_1
XANTENNA__19623__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10695_ game.CPU.applesa.ab.absxs.body_y\[87\] _04610_ _04611_ game.CPU.applesa.ab.absxs.body_y\[83\]
+ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13376__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18010_ net648 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__inv_2
X_15222_ _08787_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12434_ net1266 net377 net369 _03294_ _06310_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_340_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_340_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12365_ game.CPU.applesa.ab.absxs.body_y\[47\] net365 net362 game.CPU.applesa.ab.absxs.body_y\[44\]
+ _06241_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__o221a_1
X_15153_ net1213 net1239 game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1
+ vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__and3_1
XANTENNA__16551__X _02481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16314__B2 _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11316_ net565 _05198_ _05202_ _05204_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__o211a_1
X_14104_ net961 game.CPU.applesa.ab.check_walls.above.walls\[53\] vssd1 vssd1 vccd1
+ vccd1 _07978_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16865__A2 _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19961_ clknet_leaf_44_clk game.writer.tracker.next_frame\[556\] net1306 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[556\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19773__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15084_ net1206 net1232 game.CPU.applesa.ab.check_walls.above.walls\[112\] vssd1
+ vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__and3_1
X_12296_ _05969_ _06181_ _05971_ _05970_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14035_ net959 net798 vssd1 vssd1 vccd1 vccd1 _07909_ sky130_fd_sc_hd__xor2_1
X_18912_ clknet_leaf_3_clk _00010_ _00596_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.enable_in
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15608__A game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11247_ _03224_ net320 vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__xnor2_1
X_19892_ clknet_leaf_28_clk game.writer.tracker.next_frame\[487\] net1309 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[487\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12731__S net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14222__A2_N net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09606__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18843_ clknet_leaf_0_clk _01234_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11855__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _03300_ net538 vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__nand2_1
XANTENNA__19003__CLK net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15825__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_182_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10129_ game.CPU.randy.f1.c1.max_i\[1\] game.CPU.randy.f1.c1.count\[2\] game.CPU.randy.f1.c1.count\[1\]
+ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__o21ba_1
XANTENNA__17290__A2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12032__A game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18774_ clknet_leaf_64_clk _01191_ _00511_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[84\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12639__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13836__C1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15986_ _03420_ net442 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__nand2_1
XANTENNA__15046__C game.CPU.applesa.ab.check_walls.above.walls\[74\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13300__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17725_ game.CPU.applesa.ab.count_luck\[4\] _03091_ vssd1 vssd1 vccd1 vccd1 _03094_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14937_ _08712_ _08713_ vssd1 vssd1 vccd1 vccd1 _08714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_292_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16439__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13851__A2 _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11871__A game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17042__A2 _02670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_292_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17656_ game.CPU.kyle.L1.cnt_500hz\[9\] _03047_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14868_ game.CPU.randy.f1.c1.count\[17\] game.CPU.randy.f1.c1.count\[16\] _08653_
+ vssd1 vssd1 vccd1 vccd1 _08655_ sky130_fd_sc_hd__and3_1
XANTENNA__12686__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16607_ _02362_ _02518_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__and2b_1
X_13819_ game.writer.tracker.frame\[401\] game.writer.tracker.frame\[403\] game.writer.tracker.frame\[404\]
+ game.writer.tracker.frame\[402\] net980 net1040 vssd1 vssd1 vccd1 vccd1 _07693_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15062__B net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17587_ game.CPU.kyle.L1.cnt_20ms\[9\] game.CPU.kyle.L1.cnt_20ms\[7\] _03007_ game.CPU.kyle.L1.cnt_20ms\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__or4b_1
XFILLER_0_159_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14799_ _08612_ _08613_ vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_271_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19326_ clknet_leaf_72_clk net1426 _00931_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twomode.number\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_329_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16538_ net202 net146 _02389_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__and3_1
XANTENNA__11614__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16445__Y _02405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_311_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19257_ clknet_leaf_57_clk _01325_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.count_luck\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16469_ net2006 _02420_ _02422_ _02273_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[57\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_332_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09010_ game.CPU.applesa.ab.absxs.body_x\[109\] vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__inv_2
XANTENNA__13367__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18208_ net665 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_344_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19188_ clknet_leaf_66_clk _01306_ _00850_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.start_enable
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10934__B net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14406__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11917__A2 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18139_ net635 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold102 game.writer.tracker.frame\[202\] vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 game.writer.tracker.frame\[547\] vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold124 game.writer.tracker.frame\[354\] vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11111__A game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16856__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 game.writer.tracker.frame\[500\] vssd1 vssd1 vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12590__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold146 game.writer.tracker.frame\[370\] vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold157 game.writer.tracker.frame\[434\] vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 game.writer.tracker.frame\[495\] vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold179 game.writer.tracker.frame\[262\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09912_ net1092 net1100 net1109 _04147_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_282_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12878__A0 game.writer.tracker.frame\[48\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout604 net624 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_2
Xfanout615 net616 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_4
Xfanout626 net633 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__buf_4
XANTENNA__09516__A net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20032_ net1380 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_298_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ net1096 _03248_ _03315_ net1146 vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__o22a_1
Xfanout637 net638 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__buf_4
Xfanout648 net651 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_4
Xfanout659 net660 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_4
XANTENNA__14141__B _07953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17281__A2 _02576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ net891 game.CPU.applesa.ab.YMAX\[0\] net1171 net897 vssd1 vssd1 vccd1 vccd1
+ _04017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_280_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13980__B net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13472__S net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16349__A _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13842__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_X net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_A net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17033__A2 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10656__A2 _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12596__B net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16068__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19620__RESET_B net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_293_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16792__A1 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19646__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_X net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_235_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11005__B net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_69_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09208_ game.CPU.applesa.ab.check_walls.above.walls\[146\] vssd1 vssd1 vccd1 vccd1
+ _03457_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18670__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19796__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10480_ _04358_ _04578_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__or2_4
XANTENNA__14316__B net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09139_ game.CPU.applesa.ab.check_walls.above.walls\[18\] vssd1 vssd1 vccd1 vccd1
+ _03388_ sky130_fd_sc_hd__inv_2
XANTENNA__17908__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_301_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12150_ game.CPU.applesa.ab.check_walls.above.walls\[132\] net551 vssd1 vssd1 vccd1
+ vccd1 _06037_ sky130_fd_sc_hd__or2_1
XANTENNA__14307__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout880_X net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19026__CLK net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_X net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ game.CPU.applesa.ab.absxs.body_y\[4\] net534 vssd1 vssd1 vccd1 vccd1 _04991_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__11956__A game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12655__A2_N net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _05951_ _05952_ _05957_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_246_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11032_ _03335_ net404 vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09426__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20003__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15582__A2_N net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17272__A2 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15840_ _03386_ net271 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_290_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19176__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16480__B1 _02429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15771_ _03253_ net348 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13294__B1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12983_ net246 _06846_ _06851_ _06856_ net187 vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__a311o_2
XFILLER_0_231_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19708__RESET_B net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12097__B2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14491__C1 _08364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17510_ _04638_ _02784_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__and2b_1
XFILLER_0_262_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15163__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14722_ game.CPU.randy.counter1.count1\[6\] _08553_ vssd1 vssd1 vccd1 vccd1 _08556_
+ sky130_fd_sc_hd__or2_1
X_18490_ net588 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__inv_2
X_11934_ game.CPU.applesa.ab.check_walls.above.walls\[165\] net305 vssd1 vssd1 vccd1
+ vccd1 _05822_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_335_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _02772_ _02778_ _02817_ _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a31o_1
XFILLER_0_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14653_ _08487_ _08490_ vssd1 vssd1 vccd1 vccd1 _08492_ sky130_fd_sc_hd__nor2_1
XANTENNA__16783__A1 _02462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11865_ game.CPU.applesa.ab.check_walls.above.walls\[6\] net303 vssd1 vssd1 vccd1
+ vccd1 _05753_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16546__X _02477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_257_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13597__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13604_ _07476_ _07477_ net503 vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__mux2_1
X_10816_ _03355_ net233 vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__nor2_1
X_17372_ _02796_ _02800_ _02793_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__a21oi_1
X_14584_ game.CPU.clock1.counter\[9\] game.CPU.clock1.counter\[14\] game.CPU.clock1.counter\[16\]
+ game.CPU.clock1.counter\[21\] vssd1 vssd1 vccd1 vccd1 _08446_ sky130_fd_sc_hd__and4_1
X_11796_ net575 _05440_ _05444_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_94_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19111_ net1180 _00150_ _00782_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[156\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_55_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16323_ _02316_ net199 _01516_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13535_ net510 _07405_ _07406_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__and3_1
XFILLER_0_184_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15610__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10747_ net936 game.CPU.applesa.ab.absxs.body_y\[100\] net234 _04718_ vssd1 vssd1
+ vccd1 vccd1 _01039_ sky130_fd_sc_hd__a31o_1
XANTENNA__16535__B2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19042_ net1189 _00273_ _00713_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[87\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_313_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16254_ net1906 _02260_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[4\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13466_ _07338_ _07339_ net514 vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__mux2_1
X_10678_ _03288_ net233 vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19078__Q game.CPU.applesa.ab.check_walls.above.walls\[123\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14226__B net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15205_ game.CPU.applesa.normal1.number\[2\] _08768_ vssd1 vssd1 vccd1 vccd1 _08773_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_298_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12417_ game.CPU.applesa.ab.absxs.body_x\[32\] net381 vssd1 vssd1 vccd1 vccd1 _06294_
+ sky130_fd_sc_hd__xnor2_1
X_16185_ game.CPU.applesa.ab.check_walls.above.walls\[105\] net475 net466 game.CPU.applesa.ab.check_walls.above.walls\[106\]
+ _02157_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__o221a_1
X_13397_ net281 _07264_ _07270_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_211_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12027__A _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_301_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_346_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15136_ net1209 net1235 game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1
+ vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__and3_1
XFILLER_0_140_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12348_ game.CPU.applesa.ab.absxs.body_x\[37\] net376 vssd1 vssd1 vccd1 vccd1 _06225_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10583__A1 game.CPU.applesa.ab.absxs.body_x\[114\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19806__Q game.writer.tracker.frame\[401\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18710__Q game.CPU.applesa.ab.absxs.body_x\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19944_ clknet_leaf_38_clk game.writer.tracker.next_frame\[539\] net1329 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[539\] sky130_fd_sc_hd__dfrtp_1
X_12279_ net805 net418 vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__xnor2_1
X_15067_ net1220 net1245 game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1
+ vccd1 vccd1 _00092_ sky130_fd_sc_hd__and3_1
XANTENNA__19519__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13521__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ net881 game.CPU.applesa.ab.check_walls.above.walls\[185\] net782 net868 _07891_
+ vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__a221o_1
XANTENNA__09336__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11585__B net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15057__B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19875_ clknet_leaf_21_clk game.writer.tracker.next_frame\[470\] net1318 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[470\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17799__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11532__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_276_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17263__A2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10886__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18826_ clknet_leaf_2_clk _01217_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dfxtp_1
XANTENNA__14077__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16471__B1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18757_ clknet_leaf_53_clk _01174_ _00494_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[47\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13285__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15969_ game.CPU.applesa.ab.absxs.body_x\[66\] net468 vssd1 vssd1 vccd1 vccd1 _01981_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19669__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19190__D net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17015__A2 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17708_ _03077_ _03078_ _03079_ _03359_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__a22oi_1
XANTENNA__15073__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_357_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09490_ net892 net782 game.CPU.applesa.ab.check_walls.above.walls\[190\] net902 vssd1
+ vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__a22o_1
XANTENNA__11835__B2 game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18688_ clknet_leaf_62_clk _01105_ _00425_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_349_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09071__A game.CPU.applesa.ab.absxs.body_y\[106\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_81_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17639_ _08801_ net194 _03039_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__and3b_1
XANTENNA__16774__A1 _02435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_336_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16456__X _02413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18384__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_322_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18693__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16616__B _02370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19309_ net1164 _00033_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.out_random_2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10945__A game.CPU.applesa.ab.absxs.body_y\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout137_A _02233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19049__CLK net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_230_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1046_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13760__B2 game.writer.tracker.frame\[129\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15248__A _00293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19199__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14152__A _07799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_245_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1213_A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13512__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 net402 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_4
Xfanout412 net413 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_4
Xfanout423 net424 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_4
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_4
XANTENNA_fanout673_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 _08427_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_272_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_271_Right_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20015_ net1276 vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
X_09826_ net1159 game.CPU.applesa.ab.absxs.body_y\[12\] vssd1 vssd1 vccd1 vccd1 _04069_
+ sky130_fd_sc_hd__nand2_1
Xfanout467 net470 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__clkbuf_8
Xfanout478 net479 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_4
Xfanout489 net494 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_260_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_241_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09757_ net1086 game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1 vccd1
+ vccd1 _04000_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout461_X net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_241_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout938_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17006__A2 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_240_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09688_ net1158 game.CPU.applesa.ab.absxs.body_y\[4\] vssd1 vssd1 vccd1 vccd1 _03931_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_178_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16765__A1 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12894__X _06768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18294__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_327_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11650_ net744 _05538_ _05536_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10601_ net754 _04588_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__nor2_1
Xfanout63 net64 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_2
X_11581_ _05455_ _05456_ _05462_ _05469_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout74 net75 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16517__B2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout85 _02669_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14327__A game.CPU.applesa.ab.absxs.body_y\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_330_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout96 net97 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_2
X_13320_ net211 _07193_ _07192_ net287 vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10532_ _04358_ _04638_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__nor2_2
XFILLER_0_24_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10801__A2 _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17190__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10574__B net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13251_ game.writer.tracker.frame\[470\] game.writer.tracker.frame\[471\] net1014
+ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10463_ _03227_ _04594_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16542__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12554__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ game.CPU.applesa.ab.check_walls.above.walls\[197\] net548 vssd1 vssd1 vccd1
+ vccd1 _06088_ sky130_fd_sc_hd__xnor2_1
X_13182_ game.writer.tracker.frame\[414\] game.writer.tracker.frame\[415\] net1035
+ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__mux2_1
X_10394_ net902 game.CPU.apple_location\[6\] game.CPU.apple_location\[1\] net914 _04545_
+ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__o221a_1
XANTENNA__10565__A1 game.CPU.applesa.ab.absxs.body_x\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10565__B2 game.CPU.applesa.ab.absxs.body_x\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12133_ _06017_ _06018_ _06019_ _06012_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__o31a_1
XFILLER_0_257_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15158__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14062__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17990_ net636 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13503__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16941_ _02382_ net92 _02653_ net1504 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[298\]
+ sky130_fd_sc_hd__a22o_1
X_12064_ game.CPU.applesa.ab.check_walls.above.walls\[127\] net294 net288 net794 vssd1
+ vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__o22a_1
XANTENNA__18566__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ game.CPU.applesa.ab.absxs.body_x\[54\] net409 net546 game.CPU.applesa.ab.absxs.body_x\[55\]
+ _04904_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_166_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19660_ clknet_leaf_23_clk game.writer.tracker.next_frame\[255\] net1347 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[255\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_341_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19811__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16872_ _02549_ net108 _02629_ net1836 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[253\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_263_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout990 net992 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_4
X_18611_ clknet_leaf_63_clk _01028_ _00348_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[97\]
+ sky130_fd_sc_hd__dfrtp_4
X_15823_ _01830_ _01831_ _01832_ _01834_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__or4_1
X_19591_ clknet_leaf_36_clk game.writer.tracker.next_frame\[186\] net1355 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[186\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_216_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19542__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18542_ net611 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__inv_2
X_15754_ game.CPU.applesa.ab.check_walls.above.walls\[7\] net434 vssd1 vssd1 vccd1
+ vccd1 _01766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12966_ _06833_ _06838_ _06839_ net279 net247 vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__o221a_2
XANTENNA__19961__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16205__B1 _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14705_ game.CPU.randy.counter1.count1\[18\] net266 _08537_ _08543_ vssd1 vssd1 vccd1
+ vccd1 _08544_ sky130_fd_sc_hd__o22a_1
XFILLER_0_169_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11917_ net829 net313 net308 net830 vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__a22o_1
X_18473_ net638 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__inv_2
XFILLER_0_358_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16756__A1 _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15685_ _03224_ net349 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__xnor2_1
X_12897_ _06767_ _06769_ net689 vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17424_ _04483_ _02825_ _02833_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__and3_1
XFILLER_0_169_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14636_ game.CPU.clock1.counter\[18\] _08479_ vssd1 vssd1 vccd1 vccd1 _08480_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11848_ game.CPU.applesa.ab.check_walls.above.walls\[53\] net308 vssd1 vssd1 vccd1
+ vccd1 _05736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_200_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16436__B _02318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17355_ _04638_ _02784_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__and2_1
X_14567_ net436 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.abduyd.next_wall\[7\]
+ sky130_fd_sc_hd__clkinv_8
X_11779_ net569 _05224_ _05225_ _05228_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_119_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16306_ net1887 net720 _02304_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[12\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_190_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13518_ _07372_ _07373_ net216 vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__mux2_1
XANTENNA__13990__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17286_ net176 _02258_ net56 _02752_ net1771 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[544\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__13990__B2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17181__A1 _02483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14498_ _03209_ net1044 net868 game.CPU.apple_location\[4\] _08371_ vssd1 vssd1 vccd1
+ vccd1 _08372_ sky130_fd_sc_hd__a221o_1
XANTENNA__10484__B _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19025_ net1196 _00255_ _00696_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[70\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_298_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16237_ net507 net835 _02226_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a21oi_4
Xclkload11 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 clkload11/X sky130_fd_sc_hd__clkbuf_4
X_13449_ net704 _07031_ _07322_ net512 vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__o211a_1
Xclkload22 clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__clkinv_16
XANTENNA_max_cap357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload33 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 clkload33/X sky130_fd_sc_hd__clkbuf_4
Xclkload44 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload55 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__inv_12
XANTENNA__19341__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12545__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_298_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload66 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__clkinv_16
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16168_ _03235_ net345 net341 _03302_ _02152_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__o221a_1
XANTENNA__09410__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10556__A1 game.CPU.applesa.ab.absxs.body_x\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10556__B2 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18909__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15119_ net1207 net1230 game.CPU.applesa.ab.check_walls.above.walls\[147\] vssd1
+ vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_58_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15068__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08990_ game.CPU.applesa.ab.absxs.body_x\[61\] vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__inv_2
X_16099_ game.CPU.applesa.ab.absxs.body_x\[19\] net460 net440 game.CPU.applesa.ab.absxs.body_y\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__o22a_1
XFILLER_0_282_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_267_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14298__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19927_ clknet_leaf_48_clk game.writer.tracker.next_frame\[522\] net1301 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[522\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_239_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18379__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19491__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_317_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17236__A2 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19858_ clknet_leaf_20_clk game.writer.tracker.next_frame\[453\] net1317 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[453\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_242_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_305_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12698__Y _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16444__B1 _02404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ net927 game.CPU.applesa.ab.absxs.body_x\[119\] game.CPU.applesa.ab.absxs.body_x\[117\]
+ net917 _03850_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_143_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18809_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[12\] _00546_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19789_ clknet_leaf_24_clk game.writer.tracker.next_frame\[384\] net1345 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[384\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_222_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15798__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13353__S0 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09542_ net910 game.CPU.applesa.ab.XMAX\[0\] game.CPU.applesa.ab.XMAX\[1\] net914
+ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__a22o_1
XANTENNA__11808__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12220__A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11808__B2 game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_270_Left_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10659__B _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_203_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16747__A1 _02390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09473_ _03709_ _03712_ _03713_ _03715_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__or4_1
XANTENNA__11284__A2 _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_277_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12481__B2 game.CPU.applesa.ab.absxs.body_y\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_333_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout254_A _05207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_219_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_290_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16346__B _06573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11036__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout421_A _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout519_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload5 clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_154_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17172__A1 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10795__B2 game.CPU.applesa.ab.absxs.body_y\[38\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13986__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_340_Right_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16362__A _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1049_X net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout790_A game.CPU.applesa.ab.check_walls.above.walls\[148\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18589__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16081__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11744__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19834__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1216_X net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14143__D1 _07745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_243_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1207 net1208 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__clkbuf_2
Xfanout220 net222 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_4
Xfanout1218 game.CPU.walls.rand_wall.start_enable vssd1 vssd1 vccd1 vccd1 net1218
+ sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout231 net232 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1229 net1232 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__clkbuf_2
XANTENNA__18289__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_2
XFILLER_0_227_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17227__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout253 _05210_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_4
Xfanout264 _08810_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_245_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout275 _06610_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_2
Xfanout286 net287 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_2
XANTENNA__19984__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09704__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09809_ net924 game.CPU.applesa.ab.check_walls.above.walls\[107\] net801 net903 vssd1
+ vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__a22o_1
Xfanout297 net298 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_2
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16986__A1 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11251__A1_N game.CPU.applesa.ab.absxs.body_x\[114\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12820_ _06692_ _06693_ net511 vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_307_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09423__B game.CPU.applesa.ab.check_walls.above.walls\[112\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15144__C net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12751_ game.writer.tracker.frame\[74\] game.writer.tracker.frame\[75\] net1010 vssd1
+ vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_243_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13660__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14983__C game.CPU.applesa.ab.check_walls.above.walls\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11702_ net566 _05589_ _05588_ _05586_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__o211a_1
XANTENNA__10483__B1 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_328_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15470_ _01461_ _01496_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__nand2_1
X_12682_ net1075 net1065 vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__xor2_4
XFILLER_0_96_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_254_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14421_ game.CPU.applesa.ab.absxs.body_x\[110\] net880 net858 game.CPU.applesa.ab.absxs.body_y\[111\]
+ vssd1 vssd1 vccd1 vccd1 _08295_ sky130_fd_sc_hd__o22a_1
XFILLER_0_328_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11633_ game.CPU.applesa.ab.check_walls.above.walls\[157\] net315 vssd1 vssd1 vccd1
+ vccd1 _05522_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14057__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17140_ net185 _02410_ net80 _02714_ net1514 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[436\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__19364__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13972__A1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14352_ game.CPU.applesa.ab.absxs.body_x\[33\] net1061 vssd1 vssd1 vccd1 vccd1 _08226_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__17163__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11564_ _05450_ _05451_ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__or3_1
XANTENNA__13972__B2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10786__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13303_ _07175_ _07176_ net481 vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17071_ _02452_ net59 _02694_ net2028 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[387\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10515_ _03197_ net849 _04174_ _04609_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__o31a_1
XANTENNA__10872__X game.CPU.randy.counter1.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11495_ _05383_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14283_ game.CPU.applesa.ab.absxs.body_x\[86\] net877 net983 _03298_ vssd1 vssd1
+ vccd1 vccd1 _08157_ sky130_fd_sc_hd__a22o_1
XANTENNA__16910__A1 _02486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16272__A _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13185__C1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16022_ game.CPU.applesa.ab.absxs.body_y\[39\] net436 vssd1 vssd1 vccd1 vccd1 _02034_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13234_ _07104_ _07105_ _07106_ _07107_ net488 net686 vssd1 vssd1 vccd1 vccd1 _07108_
+ sky130_fd_sc_hd__mux4_1
X_10446_ net1123 net1124 vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__or2_2
XFILLER_0_311_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10538__A1 game.CPU.applesa.ab.absxs.body_x\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_343_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10538__B2 game.CPU.applesa.ab.absxs.body_x\[40\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13165_ _07035_ _07036_ _07038_ _07037_ net498 net690 vssd1 vssd1 vccd1 vccd1 _07039_
+ sky130_fd_sc_hd__mux4_1
X_10377_ net1153 game.CPU.apple_location2\[4\] vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__and2_1
XFILLER_0_268_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ _05990_ _05991_ _05992_ _06002_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__a31o_1
X_13096_ _06968_ _06969_ net501 vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_264_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17973_ net643 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__inv_2
XFILLER_0_209_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18199__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12024__B net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19712_ clknet_leaf_35_clk game.writer.tracker.next_frame\[307\] net1339 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[307\] sky130_fd_sc_hd__dfrtp_1
X_16924_ _02348_ _02643_ _02649_ net1949 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[285\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17218__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12047_ _05923_ _05924_ _05925_ _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__o31a_1
XFILLER_0_224_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12160__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_284_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output50_A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16855_ _02538_ net102 _02623_ game.writer.tracker.frame\[241\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[241\] sky130_fd_sc_hd__a22o_1
X_19643_ clknet_leaf_15_clk game.writer.tracker.next_frame\[238\] net1288 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[238\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15806_ game.CPU.applesa.ab.check_walls.above.walls\[63\] net434 vssd1 vssd1 vccd1
+ vccd1 _01818_ sky130_fd_sc_hd__nor2_1
X_19574_ clknet_leaf_49_clk game.writer.tracker.next_frame\[169\] net1279 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[169\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_217_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16786_ _02461_ net108 _02596_ net1777 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[199\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15054__C game.CPU.applesa.ab.check_walls.above.walls\[82\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13998_ _07866_ _07867_ _07870_ _07871_ vssd1 vssd1 vccd1 vccd1 _07872_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_179_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18525_ net583 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_354_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15737_ _03472_ net343 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16729__A1 _02512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ _06745_ _06747_ net676 vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__mux2_1
XANTENNA__11266__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16729__B2 game.writer.tracker.frame\[161\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16447__A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_319_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13570__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_72_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18456_ net654 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__inv_2
X_15668_ game.CPU.applesa.ab.check_walls.above.walls\[109\] net445 vssd1 vssd1 vccd1
+ vccd1 _01680_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19707__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14204__A2 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17407_ _02778_ _02833_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__nand2_1
X_14619_ _08469_ net741 _08468_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[11\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__15070__B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18387_ net618 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15599_ net799 net449 net465 game.CPU.applesa.ab.check_walls.above.walls\[114\] vssd1
+ vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_172_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17338_ _08908_ net576 _02765_ _02768_ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__o22a_1
XFILLER_0_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17154__A1 _02432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18731__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11103__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19857__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_287_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17269_ net183 net117 _02486_ _02748_ net1668 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[531\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_342_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16901__A1 _02237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19008_ net1194 _00236_ _00679_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[53\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_178_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10529__A1 game.CPU.applesa.ab.absxs.body_x\[53\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10529__B2 net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10942__B net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload39_A clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_307_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_302_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09508__B game.CPU.applesa.ab.absxs.body_y\[50\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_178_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16665__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_227_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18881__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08973_ game.CPU.randy.f1.state\[0\] vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__inv_2
XANTENNA__17209__A2 _02369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold17 game.CPU.down_button.eD1.Q1 vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 game.CPU.applesa.twomode.number\[4\] vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 game.CPU.applesa.normal1.number\[2\] vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_279_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09524__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16968__A1 _02432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10701__A1 game.CPU.applesa.ab.absxs.body_y\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Left_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17090__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13326__S0 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16432__A3 _02394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16628__Y _02533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09525_ net920 game.CPU.applesa.ab.check_walls.above.walls\[122\] net794 net903 _03767_
+ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__a221o_1
XANTENNA__12454__A1 game.CPU.applesa.ab.absxs.body_x\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1280_A net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_63_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout636_A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19387__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ net917 game.CPU.applesa.ab.absxs.body_x\[69\] game.CPU.applesa.ab.absxs.body_x\[70\]
+ net923 vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_80_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16076__B net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09387_ net1126 net786 vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17145__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10768__B2 game.CPU.applesa.ab.absxs.body_y\[76\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1333_X net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10300_ game.CPU.clock1.game_state\[0\] net1264 vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__and2b_1
XFILLER_0_277_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11280_ _05106_ _05107_ _05109_ _05110_ _05112_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11717__B1 game.CPU.applesa.ab.apple_possible\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14324__B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ game.CPU.applesa.ab.count_luck\[7\] game.CPU.applesa.ab.count_luck\[5\] game.CPU.applesa.ab.count_luck\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__or3b_1
XFILLER_0_293_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_292_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15139__C net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10162_ _04347_ _04352_ _04354_ _04356_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__and4_1
XFILLER_0_246_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1004 net1005 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__clkbuf_4
Xfanout1015 net1016 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_4
Xfanout1026 net1029 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13565__S0 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14978__C game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout1037 net1041 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_4
X_10093_ _04295_ _04297_ _04299_ _04300_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__and4bb_1
X_14970_ _03362_ game.CPU.walls.rand_wall.logic_enable net1243 vssd1 vssd1 vccd1 vccd1
+ _08747_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout72_X net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1048 net1049 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14340__A game.CPU.applesa.ab.absxs.body_y\[38\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1059 game.CPU.applesa.x\[2\] vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_163_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13921_ net1052 _03459_ _03461_ net958 vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__a22o_1
XANTENNA__11683__B net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16959__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_260_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16640_ net145 _02398_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852_ game.writer.tracker.frame\[562\] net842 net836 game.writer.tracker.frame\[561\]
+ net274 vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_3_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18604__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10299__B game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14994__B net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14434__A2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12803_ game.writer.tracker.frame\[370\] game.writer.tracker.frame\[371\] net1012
+ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16571_ _02243_ _02494_ net728 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__o21a_1
X_13783_ _07655_ _07656_ net498 vssd1 vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
X_10995_ game.CPU.applesa.ab.absxs.body_y\[44\] net535 vssd1 vssd1 vccd1 vccd1 _04885_
+ sky130_fd_sc_hd__or2_1
XANTENNA__13390__S net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09310__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18310_ net621 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
X_15522_ net992 net853 net699 _01542_ _01543_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__o221a_1
XANTENNA__09310__B2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12734_ net872 _06572_ net865 vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__a21oi_4
X_19290_ clknet_leaf_4_clk _01334_ _00909_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.max_i\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_44_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10586__Y _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18241_ net650 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XFILLER_0_355_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15453_ _08914_ _01476_ _01479_ _01472_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__o211a_1
XANTENNA__18754__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12665_ _06503_ _06507_ _06523_ _06541_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_100_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_343_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13945__A1 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14404_ _08269_ _08270_ _08271_ _08272_ vssd1 vssd1 vccd1 vccd1 _08278_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_174_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ net781 net259 vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__xnor2_1
X_18172_ net602 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__inv_2
XANTENNA__17136__A1 _02398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15384_ _08924_ _08925_ vssd1 vssd1 vccd1 vccd1 _08926_ sky130_fd_sc_hd__nor2_1
XANTENNA__13945__B2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12596_ game.CPU.applesa.ab.absxs.body_y\[108\] net361 vssd1 vssd1 vccd1 vccd1 _06473_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12019__B net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17123_ _02375_ net57 _02709_ net2026 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[424\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14335_ _08200_ _08201_ _08207_ _08208_ vssd1 vssd1 vccd1 vccd1 _08209_ sky130_fd_sc_hd__a211o_1
X_11547_ _05424_ _05425_ _05434_ _05435_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__or4_1
XFILLER_0_123_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15698__A1 game.CPU.applesa.ab.absxs.body_x\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17054_ _02425_ _02670_ net731 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__o21a_1
Xhold509 game.writer.tracker.frame\[132\] vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09609__A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15698__B2 game.CPU.applesa.ab.absxs.body_y\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_213_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14266_ _08137_ _08138_ _08139_ vssd1 vssd1 vccd1 vccd1 _08140_ sky130_fd_sc_hd__and3_1
X_11478_ game.CPU.applesa.ab.check_walls.above.walls\[49\] net771 vssd1 vssd1 vccd1
+ vccd1 _05367_ sky130_fd_sc_hd__xor2_1
XANTENNA__19904__RESET_B net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14234__B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__B1 _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16005_ game.CPU.applesa.ab.absxs.body_x\[60\] net271 vssd1 vssd1 vccd1 vccd1 _02017_
+ sky130_fd_sc_hd__nand2_1
X_13217_ game.writer.tracker.frame\[422\] game.writer.tracker.frame\[423\] net1024
+ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__mux2_1
X_10429_ game.CPU.right_button.eD1.Q1 _03365_ _04567_ net1078 vssd1 vssd1 vccd1 vccd1
+ _04574_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_283_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16730__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15049__C net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14197_ _08064_ _08065_ _08067_ _08068_ vssd1 vssd1 vccd1 vccd1 _08071_ sky130_fd_sc_hd__or4_1
XFILLER_0_296_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16647__B1 _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13148_ net512 _07019_ _07021_ net214 vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__o211a_1
XANTENNA__16111__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14122__A1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__A game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14122__B2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_185_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16662__A3 _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13079_ _06949_ _06950_ net678 vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17956_ net642 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12133__B1 _06012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_302_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16907_ _02479_ _02644_ net728 vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__o21a_1
XANTENNA__11593__B net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17887_ net614 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__inv_2
XANTENNA__11487__A2 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19626_ clknet_leaf_27_clk game.writer.tracker.next_frame\[221\] net1321 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[221\] sky130_fd_sc_hd__dfrtp_1
X_16838_ net1525 _02613_ _02615_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[233\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16448__Y _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_339_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16769_ _02428_ net64 _02591_ net1779 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[188\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_314_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19557_ clknet_leaf_34_clk game.writer.tracker.next_frame\[152\] net1329 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[152\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13633__A0 game.writer.tracker.frame\[49\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_177_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_200_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09310_ net899 game.CPU.applesa.ab.absxs.body_y\[53\] game.CPU.applesa.ab.absxs.body_y\[52\]
+ net893 _03546_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15081__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18508_ net579 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_274_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19488_ clknet_leaf_23_clk game.writer.tracker.next_frame\[83\] net1336 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[83\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_216_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09241_ game.CPU.walls.abc.number_out\[2\] vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__inv_2
XFILLER_0_319_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18439_ net588 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_196_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18392__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10462__A3 _04594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16905__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09172_ game.CPU.applesa.ab.check_walls.above.walls\[72\] vssd1 vssd1 vccd1 vccd1
+ _03421_ sky130_fd_sc_hd__inv_2
XANTENNA__13936__A1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17127__A1 _02299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13936__B2 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_313_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14023__A1_N net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout217_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_259_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16886__B1 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09519__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14361__A1 game.CPU.applesa.ab.absxs.body_x\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_275_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput18 net18 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XFILLER_0_339_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_285_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16640__A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1126_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_227_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout586_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14113__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__A game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13547__S0 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14113__B2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ game.CPU.apple_location2\[1\] vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__inv_2
XANTENNA__18627__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12124__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17063__B1 _02689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09541__X _03784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11008__B net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15703__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout920_A net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18777__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_296_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09508_ net1142 game.CPU.applesa.ab.absxs.body_y\[50\] vssd1 vssd1 vccd1 vccd1 _03751_
+ sky130_fd_sc_hd__or2_1
X_10780_ game.CPU.applesa.ab.absxs.body_y\[58\] net327 _04721_ net933 vssd1 vssd1
+ vccd1 vccd1 _01009_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_238_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_344_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09439_ net1112 game.CPU.applesa.ab.absxs.body_x\[56\] vssd1 vssd1 vccd1 vccd1 _03682_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_240_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12450_ game.CPU.applesa.ab.absxs.body_x\[48\] net384 vssd1 vssd1 vccd1 vccd1 _06327_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__17118__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16534__B _02300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11401_ net567 _05282_ _05288_ _05289_ _05285_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a221o_1
X_12381_ _06252_ _06257_ _06253_ _06255_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__or4b_1
XANTENNA__11402__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14120_ _07988_ _07992_ _07993_ vssd1 vssd1 vccd1 vccd1 _07994_ sky130_fd_sc_hd__or3_1
XFILLER_0_151_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11332_ net810 net249 vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__nor2_1
XANTENNA__11678__B net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_327_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14054__B net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19402__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14051_ net868 game.CPU.applesa.ab.check_walls.above.walls\[196\] net780 net857 vssd1
+ vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__a22o_1
XANTENNA__15718__X _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11263_ game.CPU.applesa.ab.absxs.body_y\[103\] net397 _04819_ game.CPU.applesa.ab.absxs.body_y\[100\]
+ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_265_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_249_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16550__A net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12363__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ game.writer.tracker.frame\[542\] game.writer.tracker.frame\[543\] net1021
+ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_249_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16629__B1 _02533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10214_ _04376_ _04378_ _04377_ _04373_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__a211o_1
X_11194_ _05080_ _05083_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_42_Left_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13385__S net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11694__A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17810_ _08884_ _03144_ _08898_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__o21ba_1
X_10145_ game.CPU.randy.f1.c1.count\[9\] game.CPU.randy.f1.c1.count\[8\] _04326_ _04339_
+ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__or4_2
X_18790_ clknet_leaf_9_clk _01205_ _00527_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_219_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14070__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19552__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_265_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17741_ net1955 _03099_ _03104_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09164__A net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ _04272_ _04278_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__xor2_1
X_14953_ game.CPU.walls.rand_wall.count_luck\[4\] game.CPU.walls.rand_wall.count_luck\[3\]
+ vssd1 vssd1 vccd1 vccd1 _08730_ sky130_fd_sc_hd__nand2_1
XANTENNA__11469__A2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16549__X _02479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13863__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17054__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13904_ net958 net795 vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_50_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17672_ _03488_ _04255_ _08695_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__or3_1
X_14884_ net1134 _08428_ vssd1 vssd1 vccd1 vccd1 _08661_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16268__Y _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09451__X _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15604__A1 game.CPU.applesa.ab.check_walls.above.walls\[115\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16623_ net199 _02528_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__nand2_1
X_19411_ clknet_leaf_48_clk game.writer.tracker.next_frame\[6\] net1295 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_214_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_338_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13835_ net484 _07702_ _07703_ _07704_ net279 vssd1 vssd1 vccd1 vccd1 _07709_ sky130_fd_sc_hd__a221o_1
XFILLER_0_214_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15613__B net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_281_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10429__B1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16554_ game.writer.tracker.frame\[81\] _02481_ _02483_ net129 vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[81\] sky130_fd_sc_hd__a22o_1
XANTENNA__13710__S0 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19342_ clknet_leaf_72_clk _01357_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.count\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13766_ game.writer.tracker.frame\[190\] net844 net711 game.writer.tracker.frame\[191\]
+ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__o22a_1
XFILLER_0_186_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ game.CPU.applesa.ab.absxs.body_x\[74\] net410 vssd1 vssd1 vccd1 vccd1 _04868_
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_51_Left_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14229__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_328_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15505_ net872 _01527_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__nor2_1
X_12717_ _06578_ _06590_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__xnor2_1
X_19273_ clknet_leaf_7_clk _00043_ _00903_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_16485_ _02274_ _02432_ net736 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__o21a_1
X_13697_ game.writer.tracker.frame\[473\] game.writer.tracker.frame\[475\] game.writer.tracker.frame\[476\]
+ game.writer.tracker.frame\[474\] net975 net1017 vssd1 vssd1 vccd1 vccd1 _07571_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13379__C1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18224_ net649 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__inv_2
X_15436_ _01459_ _01463_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17109__A1 _02577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12648_ game.CPU.applesa.ab.absxs.body_x\[94\] net370 game.CPU.applesa.twoapples.absxs.next_head\[6\]
+ _03296_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__a22o_1
XFILLER_0_316_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09598__A1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18155_ net635 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__inv_2
XANTENNA__09598__B2 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12456__A1_N net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18713__Q game.CPU.applesa.ab.absxs.body_x\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15367_ game.writer.updater.commands.cmd_num\[3\] _08877_ vssd1 vssd1 vccd1 vccd1
+ _08909_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12579_ game.CPU.applesa.ab.absxs.body_x\[20\] net385 vssd1 vssd1 vccd1 vccd1 _06456_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__12317__X _06203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14245__A game.CPU.applesa.ab.absxs.body_x\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_300_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17106_ _02576_ net81 _02704_ net1950 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[412\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14318_ game.CPU.applesa.ab.absxs.body_x\[59\] net874 net964 _03339_ vssd1 vssd1
+ vccd1 vccd1 _08192_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_349_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18086_ net639 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__inv_2
X_15298_ game.CPU.applesa.twomode.number\[5\] _08842_ net757 vssd1 vssd1 vccd1 vccd1
+ _08847_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold306 game.CPU.randy.f1.c1.count\[7\] vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 game.writer.tracker.frame\[60\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19082__CLK net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold328 game.writer.tracker.frame\[390\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_257_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold339 game.writer.tracker.frame\[177\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_257_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17037_ _02389_ _02516_ net119 _02682_ net1593 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[365\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__13777__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14249_ game.CPU.applesa.ab.absxs.body_x\[21\] net1063 vssd1 vssd1 vccd1 vccd1 _08123_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_309_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout808 game.CPU.applesa.ab.check_walls.above.walls\[87\] vssd1 vssd1 vccd1 vccd1
+ net808 sky130_fd_sc_hd__clkbuf_4
Xfanout819 game.CPU.applesa.ab.check_walls.above.walls\[54\] vssd1 vssd1 vccd1 vccd1
+ net819 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13295__S net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19193__D net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13529__S0 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15076__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09770__A1 net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09790_ net1151 game.CPU.applesa.ab.absxs.body_y\[41\] vssd1 vssd1 vccd1 vccd1 _04033_
+ sky130_fd_sc_hd__xnor2_1
X_18988_ net1197 _00214_ _00659_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[33\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_252_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09074__A game.CPU.applesa.ab.absxs.body_y\[113\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_264_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_183_Right_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17939_ net657 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__inv_2
XANTENNA__16459__X _02416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13854__B1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12212__B net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18387__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16399__A2 _02370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_222_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19609_ clknet_leaf_18_clk game.writer.tracker.next_frame\[204\] net1310 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[204\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13606__A0 game.writer.tracker.frame\[289\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_198_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09802__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15523__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11880__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout167_A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13701__S0 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13082__A1 game.writer.tracker.frame\[209\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__B game.CPU.applesa.ab.check_walls.above.walls\[120\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_326_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16635__A net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19897__RESET_B net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1076_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09224_ game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1 vccd1 vccd1
+ _03473_ sky130_fd_sc_hd__inv_2
XANTENNA__13909__A1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13909__B2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_334_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16571__A2 _02494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19826__RESET_B net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_350_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09589__A1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18623__Q game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19425__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ net821 vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__inv_2
XANTENNA__09589__B2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout501_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout122_X net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14155__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1243_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_233_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12593__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09086_ game.CPU.applesa.ab.absxs.body_y\[65\] vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__inv_2
XANTENNA__13994__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16874__A3 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1129_X net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19575__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19454__Q game.writer.tracker.frame\[49\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout870_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17284__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout968_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16087__B2 game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09761__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09761__B2 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ game.CPU.apple_location2\[3\] _04208_ _04209_ net1475 vssd1 vssd1 vccd1 vccd1
+ _01376_ sky130_fd_sc_hd__a22o_1
XANTENNA__10371__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18297__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09513__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15714__A game.CPU.applesa.ab.absxs.body_y\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09513__B2 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ game.CPU.applesa.ab.check_walls.above.walls\[116\] net390 _05837_ _05305_
+ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__o211a_1
X_10901_ game.CPU.applesa.ab.check_walls.collision_right _04801_ vssd1 vssd1 vccd1
+ vccd1 _04803_ sky130_fd_sc_hd__or2_1
XFILLER_0_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11881_ net791 net299 _05761_ _05762_ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__o2111a_2
XANTENNA_fanout923_X net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13620_ _07492_ _07493_ net512 vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_315_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10832_ game.writer.control.current\[0\] game.writer.control.current\[1\] _04737_
+ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__nand3_2
XANTENNA__15152__C game.CPU.applesa.ab.check_walls.above.walls\[180\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13551_ game.writer.tracker.frame\[105\] game.writer.tracker.frame\[107\] game.writer.tracker.frame\[108\]
+ game.writer.tracker.frame\[106\] net967 net989 vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10763_ game.CPU.applesa.ab.absxs.body_y\[89\] _04590_ net329 game.CPU.applesa.ab.absxs.body_y\[85\]
+ vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_251_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12502_ game.CPU.applesa.ab.absxs.body_x\[60\] net383 vssd1 vssd1 vccd1 vccd1 _06379_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_183_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16270_ net162 _02271_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_333_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13482_ net694 _07150_ _07354_ _07355_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__a22o_1
XANTENNA__16562__A2 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19567__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ game.CPU.applesa.ab.absxs.body_y\[92\] _04601_ _04709_ game.CPU.applesa.ab.absxs.body_y\[88\]
+ vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_171_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15221_ game.CPU.applesa.normal1.counter _08783_ _08784_ _08785_ _08786_ vssd1 vssd1
+ vccd1 vccd1 _08787_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11689__A net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12433_ game.CPU.applesa.ab.absxs.body_y\[101\] net526 net360 game.CPU.applesa.ab.absxs.body_y\[100\]
+ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_341_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14065__A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12584__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15152_ net1210 net1236 game.CPU.applesa.ab.check_walls.above.walls\[180\] vssd1
+ vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__and3_1
XANTENNA__09159__A game.CPU.applesa.ab.check_walls.above.walls\[51\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_340_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19918__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12364_ game.CPU.applesa.ab.absxs.body_y\[45\] net524 game.CPU.applesa.twoapples.absxs.next_head\[4\]
+ _03311_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_285_Right_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14103_ net951 net819 vssd1 vssd1 vccd1 vccd1 _07977_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_239_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11315_ net744 _05197_ _05201_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11201__B net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19960_ clknet_leaf_44_clk game.writer.tracker.next_frame\[555\] net1306 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[555\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15522__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10880__X _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15083_ net1212 net1238 net800 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__and3_1
XANTENNA__16865__A3 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12295_ game.CPU.applesa.ab.check_walls.above.walls\[21\] net550 vssd1 vssd1 vccd1
+ vccd1 _06181_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08998__A game.CPU.applesa.ab.absxs.body_x\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14034_ net1071 game.CPU.applesa.ab.check_walls.above.walls\[112\] vssd1 vssd1 vccd1
+ vccd1 _07908_ sky130_fd_sc_hd__xnor2_1
X_18911_ clknet_leaf_3_clk _00009_ _00595_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.enable_in
+ sky130_fd_sc_hd__dfrtp_4
X_11246_ game.CPU.applesa.ab.absxs.body_x\[7\] net544 net538 game.CPU.applesa.ab.absxs.body_y\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__o22a_1
X_19891_ clknet_leaf_28_clk game.writer.tracker.next_frame\[486\] net1309 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[486\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15608__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18842_ clknet_leaf_0_clk _01233_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_276_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11177_ game.CPU.applesa.ab.absxs.body_y\[78\] net402 vssd1 vssd1 vccd1 vccd1 _05067_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10128_ game.CPU.randy.f1.c1.count\[14\] game.CPU.randy.f1.c1.count\[17\] game.CPU.randy.f1.c1.count\[16\]
+ game.CPU.randy.f1.c1.count\[18\] vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__or4_1
XANTENNA__12639__A1 game.CPU.applesa.ab.absxs.body_x\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17290__A3 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15985_ game.CPU.applesa.ab.check_walls.above.walls\[70\] net334 vssd1 vssd1 vccd1
+ vccd1 _01997_ sky130_fd_sc_hd__nand2_1
X_18773_ clknet_leaf_59_clk _01190_ _00510_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[79\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_209_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10104__Y _04311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12032__B net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12639__B2 game.CPU.applesa.ab.absxs.body_y\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09504__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14936_ _08673_ _08675_ vssd1 vssd1 vccd1 vccd1 _08713_ sky130_fd_sc_hd__xor2_1
X_10059_ net1096 _04210_ _04213_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__o21a_1
X_17724_ game.CPU.applesa.ab.count_luck\[4\] game.CPU.applesa.ab.count_luck\[3\] _03089_
+ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__and3_1
XFILLER_0_292_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11871__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17655_ game.CPU.kyle.L1.cnt_500hz\[9\] _03047_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_19_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14867_ net1551 _08653_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[16\]
+ sky130_fd_sc_hd__xor2_1
XANTENNA__15589__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13818_ game.writer.tracker.frame\[405\] game.writer.tracker.frame\[407\] game.writer.tracker.frame\[408\]
+ game.writer.tracker.frame\[406\] net981 net1037 vssd1 vssd1 vccd1 vccd1 _07692_
+ sky130_fd_sc_hd__mux4_1
X_16606_ _02236_ _02517_ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__nor2_4
XFILLER_0_225_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17586_ game.CPU.kyle.L1.cnt_20ms\[12\] _03006_ game.CPU.kyle.L1.cnt_20ms\[10\] _03005_
+ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__or4b_1
XFILLER_0_348_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14798_ game.CPU.randy.counter1.count\[7\] _08610_ net139 vssd1 vssd1 vccd1 vccd1
+ _08613_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_308_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16537_ net1755 _02469_ _02471_ net124 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[76\]
+ sky130_fd_sc_hd__a22o_1
X_19325_ clknet_leaf_72_clk _00030_ _00930_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twomode.number\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_106_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_271_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19448__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ _07621_ _07622_ net482 vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__mux2_1
XANTENNA__11614__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_319_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16468_ net172 _02421_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_193_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19256_ clknet_leaf_66_clk _01324_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.count_luck\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17750__A1 net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_332_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_289_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15419_ _08880_ _01446_ _01438_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__o21ai_1
X_18207_ net666 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_310_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19187_ net1179 _00292_ _00849_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.logic_enable
+ sky130_fd_sc_hd__dfstp_4
X_16399_ _02274_ _02370_ net721 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__o21a_1
XANTENNA__12047__X _05934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19598__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09069__A game.CPU.applesa.ab.absxs.body_y\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18138_ net631 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__inv_2
XANTENNA__09430__A1_N net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold103 game.writer.tracker.frame\[230\] vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_331_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold114 game.writer.tracker.frame\[204\] vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_252_Right_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11111__B net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_269_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold125 game.CPU.clock1.counter\[21\] vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
X_18069_ net648 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__inv_2
Xhold136 game.writer.tracker.frame\[245\] vssd1 vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12922__S net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_7_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
Xhold147 game.writer.tracker.frame\[431\] vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 game.writer.tracker.frame\[88\] vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13524__C1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09911_ net1261 game.CPU.bodymain1.Direction\[0\] vssd1 vssd1 vccd1 vccd1 _04153_
+ sky130_fd_sc_hd__nand2_1
Xhold169 game.writer.tracker.frame\[332\] vssd1 vssd1 vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_282_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12878__A1 game.writer.tracker.frame\[49\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout605 net607 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__buf_4
Xfanout616 net619 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_4
X_20031_ net1278 vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
X_09842_ _04081_ _04084_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__nand2_2
Xfanout627 net633 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__buf_2
Xfanout638 net640 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_4
Xfanout649 net650 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_4
XFILLER_0_225_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14141__C _07973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ _04008_ _04009_ _04013_ _04015_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_146_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13827__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout284_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13753__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09532__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18618__Q game.CPU.applesa.ab.absxs.body_y\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout451_A _08425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1193_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout549_A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_293_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16792__A2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12802__A1 game.writer.tracker.frame\[375\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_235_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout716_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1079_X net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16084__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09207_ game.CPU.applesa.ab.check_walls.above.walls\[144\] vssd1 vssd1 vccd1 vccd1
+ _03456_ sky130_fd_sc_hd__inv_2
XFILLER_0_323_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16652__X _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12566__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13763__C1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09138_ game.CPU.applesa.ab.check_walls.above.walls\[17\] vssd1 vssd1 vccd1 vccd1
+ _03387_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10041__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_288_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10041__B2 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11021__B net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09069_ game.CPU.applesa.ab.absxs.body_y\[15\] vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__inv_2
XANTENNA__15709__A game.CPU.applesa.ab.absxs.body_y\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11100_ game.CPU.applesa.ab.absxs.body_y\[56\] net536 vssd1 vssd1 vccd1 vccd1 _04990_
+ sky130_fd_sc_hd__or2_1
XANTENNA__15428__B _01454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _05963_ _05964_ _05965_ _05966_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__and4b_1
XANTENNA__11956__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 game.writer.tracker.frame\[63\] vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_246_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09734__A1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11031_ game.CPU.applesa.ab.absxs.body_y\[64\] net535 vssd1 vssd1 vccd1 vccd1 _04921_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__17924__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09426__B net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09734__B2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15147__C game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17272__A3 _02328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13663__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14986__C game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16480__B2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15770_ game.CPU.applesa.ab.absxs.body_y\[106\] net441 vssd1 vssd1 vccd1 vccd1 _01782_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13294__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ _06852_ _06853_ _06854_ _06855_ net238 vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__o221a_1
XANTENNA__09442__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14721_ game.CPU.randy.counter1.count1\[6\] _08553_ vssd1 vssd1 vccd1 vccd1 _08555_
+ sky130_fd_sc_hd__and2_1
X_11933_ game.CPU.applesa.ab.check_walls.above.walls\[164\] net391 vssd1 vssd1 vccd1
+ vccd1 _05821_ sky130_fd_sc_hd__xor2_1
XFILLER_0_262_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_335_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17440_ _02782_ _02839_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__and2_1
XFILLER_0_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14652_ _04351_ _08487_ vssd1 vssd1 vccd1 vccd1 _08491_ sky130_fd_sc_hd__nor2_2
XANTENNA__13046__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _05732_ _05734_ _05740_ _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__a31o_1
XANTENNA__16783__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_257_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ game.writer.tracker.frame\[269\] game.writer.tracker.frame\[271\] game.writer.tracker.frame\[272\]
+ game.writer.tracker.frame\[270\] net967 net996 vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__mux4_1
XANTENNA__11057__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_354_Right_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10815_ net936 game.CPU.applesa.ab.absxs.body_y\[113\] net233 _04731_ vssd1 vssd1
+ vccd1 vccd1 _00984_ sky130_fd_sc_hd__a31o_1
X_17371_ _02800_ _02793_ _02796_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__mux2_1
XANTENNA__13899__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14583_ game.CPU.clock1.counter\[15\] game.CPU.clock1.counter\[19\] _03521_ _08444_
+ vssd1 vssd1 vccd1 vccd1 _08445_ sky130_fd_sc_hd__or4b_1
XANTENNA__16275__A _06573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11795_ net749 _05441_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__nand2_1
X_16322_ _06571_ net842 _06607_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19110_ net1180 _00149_ _00781_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[155\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13534_ game.writer.tracker.frame\[122\] net843 net837 game.writer.tracker.frame\[121\]
+ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10746_ _03321_ net234 vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__nor2_1
XANTENNA__19740__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_314_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10280__A1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19041_ net1189 _00272_ _00712_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16253_ net1854 _02260_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[3\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_353_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13465_ _07095_ _07097_ net705 vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10677_ net935 game.CPU.applesa.ab.absxs.body_x\[113\] _04701_ _04705_ vssd1 vssd1
+ vccd1 vccd1 _01096_ sky130_fd_sc_hd__a31o_1
XFILLER_0_125_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15204_ _08772_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__inv_2
XANTENNA__12557__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12416_ _03275_ game.CPU.applesa.twoapples.absxs.next_head\[2\] vssd1 vssd1 vccd1
+ vccd1 _06293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16184_ _02133_ _02190_ _02192_ _02195_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__o211a_1
XANTENNA__12021__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13396_ net225 _07265_ _07269_ net274 vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__o211a_1
XANTENNA__12027__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15135_ net1209 net1233 game.CPU.applesa.ab.check_walls.above.walls\[163\] vssd1
+ vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__and3_1
XANTENNA__17496__B1 net1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_346_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12347_ game.CPU.applesa.ab.absxs.body_x\[39\] net529 net527 game.CPU.applesa.ab.absxs.body_y\[37\]
+ _06223_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__o221a_1
XFILLER_0_279_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19890__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10583__A2 _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13506__C1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19943_ clknet_leaf_38_clk game.writer.tracker.next_frame\[538\] net1324 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[538\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_268_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09617__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15066_ net1217 net1244 game.CPU.applesa.ab.check_walls.above.walls\[94\] vssd1 vssd1
+ vccd1 vccd1 _00091_ sky130_fd_sc_hd__and3_1
X_12278_ net806 net548 vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_130_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_266_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17248__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__A1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14017_ net1053 game.CPU.applesa.ab.check_walls.above.walls\[186\] vssd1 vssd1 vccd1
+ vccd1 _07891_ sky130_fd_sc_hd__xor2_1
X_11229_ _05115_ _05116_ _05117_ _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__a22o_1
XANTENNA__09725__B2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19874_ clknet_leaf_21_clk game.writer.tracker.next_frame\[469\] net1316 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[469\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18825_ clknet_leaf_1_clk _01216_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__dfxtp_1
XANTENNA__17263__A3 _02393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16471__B2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_269_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18756_ clknet_leaf_53_clk _01173_ _00493_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[46\]
+ sky130_fd_sc_hd__dfrtp_4
X_15968_ _03334_ net442 vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_11_clk_X clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14482__B1 _08129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17707_ _03079_ _03080_ _03082_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__and3_1
XANTENNA__15073__B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14919_ _08672_ _08674_ _08676_ _08671_ vssd1 vssd1 vccd1 vccd1 _08696_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_357_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18687_ clknet_leaf_62_clk _01104_ _00424_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__19270__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15899_ game.CPU.applesa.ab.absxs.body_y\[40\] net341 vssd1 vssd1 vccd1 vccd1 _01911_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_187_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17638_ game.CPU.kyle.L1.cnt_500hz\[0\] game.CPU.kyle.L1.cnt_500hz\[1\] game.CPU.kyle.L1.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16774__A2 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_322_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_26_clk_X clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11106__B net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_321_Right_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12917__S net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17569_ net1477 _08808_ _02993_ _00293_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__o211a_1
XFILLER_0_175_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19308_ net1165 _00032_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.out_random_2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10945__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14417__B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload69_A clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_305_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14537__B2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15734__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19239_ clknet_leaf_17_clk _00070_ _00877_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_61_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16472__X _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12218__A game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11122__A game.CPU.applesa.ab.absxs.body_y\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13745__C1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_230_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09964__A1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15529__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13760__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09527__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11776__B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_A _06596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 net403 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_2
XFILLER_0_285_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout413 net414 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_4
XFILLER_0_347_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout424 _04781_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1206_A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_8
X_20014_ net1276 vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
Xfanout446 net448 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_8
X_09825_ net1085 game.CPU.applesa.ab.absxs.body_x\[15\] vssd1 vssd1 vccd1 vccd1 _04068_
+ sky130_fd_sc_hd__xor2_1
Xfanout457 net459 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_4
XANTENNA_input4_A gpio_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout468 net470 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_4
Xfanout479 net480 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout666_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19613__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout287_X net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ _03995_ _03996_ _03997_ _03998_ _03994_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__a221o_1
XFILLER_0_241_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14473__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_241_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_240_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09687_ net1159 _03295_ _03926_ _03929_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__a211o_1
XANTENNA__12400__B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16765__A2 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19841__RESET_B net1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19763__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16366__Y _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15711__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ _04671_ game.CPU.applesa.ab.absxs.body_x\[96\] _04667_ vssd1 vssd1 vccd1
+ vccd1 _01139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout53 _02386_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_4
X_11580_ net793 net249 _05467_ _05468_ _05463_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__a221o_1
Xfanout64 net65 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12882__S0 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout75 net76 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__buf_2
XANTENNA__14327__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout86 _02638_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_4
XFILLER_0_335_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_330_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout97 _02635_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__buf_2
X_10531_ _04176_ _04627_ _04578_ _04618_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__or4b_4
XFILLER_0_134_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12128__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17190__A2 _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12539__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13250_ game.writer.tracker.frame\[466\] game.writer.tracker.frame\[467\] net1011
+ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10462_ net931 game.CPU.applesa.ab.absxs.body_x\[99\] _04594_ _04596_ vssd1 vssd1
+ vccd1 vccd1 _01202_ sky130_fd_sc_hd__a31o_1
XANTENNA__16542__B net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12201_ game.CPU.applesa.ab.check_walls.above.walls\[199\] net424 vssd1 vssd1 vccd1
+ vccd1 _06087_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ game.writer.tracker.frame\[410\] game.writer.tracker.frame\[411\] net1036
+ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__mux2_1
X_10393_ net1105 _03211_ _04543_ _04544_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__o211a_1
XANTENNA__10565__A2 _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19143__CLK net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_276_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09437__A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11762__B2 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12132_ net831 net297 net291 game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1
+ vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a22o_1
XANTENNA__15158__B net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16150__B1 _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_257_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09707__A1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16940_ _02378_ net87 _02653_ net1646 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[297\]
+ sky130_fd_sc_hd__a22o_1
X_12063_ _05947_ _05949_ _05918_ _05934_ _05942_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_257_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12711__B1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14997__B net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ game.CPU.applesa.ab.absxs.body_x\[54\] net409 _03241_ net324 vssd1 vssd1
+ vccd1 vccd1 _04904_ sky130_fd_sc_hd__a2bb2o_1
X_16871_ net152 _02428_ net107 _02629_ net1704 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[252\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_341_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19293__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout980 net981 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__buf_4
X_18610_ clknet_leaf_70_clk _01027_ _00347_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[96\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout991 net992 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15822_ net1268 net457 net449 game.CPU.applesa.ab.absxs.body_y\[88\] _01833_ vssd1
+ vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__a221o_1
X_19590_ clknet_leaf_36_clk game.writer.tracker.next_frame\[185\] net1354 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[185\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_231_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19929__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15753_ _03381_ game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 _01765_ sky130_fd_sc_hd__nor2_1
X_18541_ net612 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__inv_2
X_12965_ _06766_ _06773_ net217 vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__mux2_1
XANTENNA__12310__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11916_ game.CPU.applesa.ab.check_walls.above.walls\[12\] net393 _05802_ _05803_
+ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__a211o_1
X_14704_ _08533_ _08542_ vssd1 vssd1 vccd1 vccd1 _08543_ sky130_fd_sc_hd__nor2_1
X_15684_ _03223_ net345 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__xnor2_1
X_18472_ net637 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__inv_2
X_12896_ game.writer.tracker.frame\[30\] game.writer.tracker.frame\[31\] net1025 vssd1
+ vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14216__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09891__B1 _04064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16756__A2 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _08479_ net267 _08478_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[17\]
+ sky130_fd_sc_hd__and3b_1
X_17423_ _04483_ _02851_ _02852_ net1274 vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__a22o_1
XANTENNA__15621__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11847_ game.CPU.applesa.ab.check_walls.above.walls\[53\] net308 vssd1 vssd1 vccd1
+ vccd1 _05735_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_177_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _03488_ _04256_ _08430_ vssd1 vssd1 vccd1 vccd1 _08431_ sky130_fd_sc_hd__or3_1
X_17354_ _02773_ _02783_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__nor2_2
X_11778_ net749 _05226_ _05224_ net569 vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_119_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13517_ net241 _07357_ _07362_ _07388_ _07390_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__a32o_1
X_16305_ _02274_ _02303_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_190_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17285_ net117 net160 _02434_ _02752_ net1682 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[543\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10729_ game.CPU.applesa.ab.absxs.body_y\[30\] net330 _04714_ game.CPU.applesa.ab.absxs.body_y\[26\]
+ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__a22o_1
X_14497_ _03211_ net1069 net1060 _03210_ vssd1 vssd1 vccd1 vccd1 _08371_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16236_ net502 net836 vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__nand2_1
X_19024_ net1199 _00253_ _00695_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[69\]
+ sky130_fd_sc_hd__dfrtp_1
X_13448_ net684 _07034_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__or2_1
Xclkload12 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__inv_6
XFILLER_0_152_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload23 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__inv_8
XFILLER_0_298_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10005__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload34 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 clkload34/Y sky130_fd_sc_hd__inv_8
Xclkload45 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__bufinv_16
Xclkload56 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__inv_8
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16167_ game.CPU.applesa.ab.absxs.body_y\[76\] net449 game.CPU.walls.rand_wall.abduyd.next_wall\[7\]
+ _03299_ _02156_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__o221a_1
XFILLER_0_298_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13379_ net188 _07189_ _07229_ _07252_ net180 vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__o221a_1
Xclkload67 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__inv_8
XANTENNA__12325__X _06209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14253__A game.CPU.applesa.ab.absxs.body_y\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_140_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11753__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15118_ net1208 net1233 game.CPU.applesa.ab.check_walls.above.walls\[146\] vssd1
+ vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11596__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_53_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09347__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15068__B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16098_ game.CPU.applesa.ab.absxs.body_x\[19\] net460 net440 game.CPU.applesa.ab.absxs.body_y\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__a22o_1
XFILLER_0_267_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19636__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16692__A1 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19926_ clknet_leaf_48_clk game.writer.tracker.next_frame\[521\] net1301 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[521\] sky130_fd_sc_hd__dfrtp_1
X_15049_ net1214 net1240 net813 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_114_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11505__A1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17236__A3 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_317_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19857_ clknet_leaf_20_clk game.writer.tracker.next_frame\[452\] net1315 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[452\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_305_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_282_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09610_ net1132 game.CPU.applesa.ab.absxs.body_y\[119\] vssd1 vssd1 vccd1 vccd1 _03853_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__15084__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16444__B2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18808_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[11\] _00545_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[11\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19788_ clknet_leaf_24_clk game.writer.tracker.next_frame\[383\] net1346 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[383\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19786__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18660__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09082__A game.CPU.applesa.ab.absxs.body_y\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_20049__1368 vssd1 vssd1 vccd1 vccd1 _20049__1368/HI net1368 sky130_fd_sc_hd__conb_1
XFILLER_0_222_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09541_ _03775_ _03776_ _03778_ _03783_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__or4_2
XANTENNA__13353__S1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18739_ clknet_leaf_9_clk _01156_ _00476_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11808__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18395__A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12220__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_250_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_203_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10021__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09472_ net924 game.CPU.applesa.ab.absxs.body_x\[95\] game.CPU.applesa.ab.absxs.body_y\[93\]
+ net898 _03714_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_69_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_277_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12481__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__A3 _05164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19016__CLK net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_290_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout247_A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16346__C _06607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload6 clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__inv_12
XFILLER_0_289_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17172__A2 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1156_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10795__A2 _04690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16362__B _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13733__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Left_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18631__Q game.CPU.applesa.ab.absxs.body_y\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout202_X net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1323_A net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11744__A1 game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_288_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16132__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16683__A1 _02252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_285_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout210 net211 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_243_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1111_X net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1208 net1209 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__clkbuf_2
Xfanout221 net222 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_4
Xfanout1219 net1220 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__clkbuf_2
Xfanout232 _06591_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1209_X net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17227__A3 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout243 _06619_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15706__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout254 _05207_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_4
XANTENNA_fanout950_A game.CPU.applesa.y\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_2
XANTENNA__16435__A1 game.writer.tracker.frame\[48\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 _06610_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16435__B2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout287 _06609_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_4
XANTENNA__17632__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ net918 game.CPU.applesa.ab.check_walls.above.walls\[105\] _03439_ net1136
+ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09704__B game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 _05858_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout62_A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16986__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09739_ net1103 game.CPU.applesa.ab.check_walls.above.walls\[65\] vssd1 vssd1 vccd1
+ vccd1 _03982_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_98_Left_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_307_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_X clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12750_ game.writer.tracker.frame\[78\] game.writer.tracker.frame\[79\] net999 vssd1
+ vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__mux2_1
XANTENNA__16199__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16738__A2 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11701_ net742 _05587_ _05589_ net566 vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__a22oi_1
XANTENNA__09720__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12681_ net888 net883 vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__nor2_1
XFILLER_0_328_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_254_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ net853 game.CPU.applesa.ab.absxs.body_y\[110\] _03257_ net1050 vssd1 vssd1
+ vccd1 vccd1 _08294_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_323_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11632_ net788 net258 vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19509__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16824__Y _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14057__B game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14351_ game.CPU.applesa.ab.absxs.body_y\[34\] net949 vssd1 vssd1 vccd1 vccd1 _08225_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11563_ net780 net259 net255 game.CPU.applesa.ab.check_walls.above.walls\[198\] vssd1
+ vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13972__A2 game.CPU.applesa.ab.check_walls.above.walls\[80\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17163__A2 _02454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16553__A _02318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13302_ _06747_ _06768_ net676 vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__mux2_1
XANTENNA__10786__A2 game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17070_ _02444_ net60 net559 vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a21oi_2
X_10514_ net1078 _03527_ _04628_ _04156_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__o31a_1
X_14282_ game.CPU.applesa.ab.absxs.body_y\[86\] net947 vssd1 vssd1 vccd1 vccd1 _08156_
+ sky130_fd_sc_hd__or2_1
X_11494_ game.CPU.applesa.ab.check_walls.above.walls\[168\] net776 vssd1 vssd1 vccd1
+ vccd1 _05383_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_311_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16272__B net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13388__S net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19286__D net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16021_ _03245_ net352 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19659__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ game.writer.tracker.frame\[506\] game.writer.tracker.frame\[507\] net1030
+ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__mux2_1
XANTENNA__15169__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09928__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_268_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10445_ net1123 game.CPU.bodymain1.main.score\[0\] vssd1 vssd1 vccd1 vccd1 _04580_
+ sky130_fd_sc_hd__nor2_2
XANTENNA__12932__A0 _06710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10538__A2 _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_343_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09167__A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13164_ game.writer.tracker.frame\[190\] game.writer.tracker.frame\[191\] net1038
+ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__mux2_1
XANTENNA__16123__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10376_ net906 game.CPU.apple_location2\[7\] game.CPU.apple_location2\[5\] net897
+ _04527_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__o221a_1
XANTENNA__12305__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ _06001_ _05994_ _05993_ _05995_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_265_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13095_ _06965_ _06967_ net693 vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__mux2_1
X_17972_ net663 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_207_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18683__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19711_ clknet_leaf_35_clk game.writer.tracker.next_frame\[306\] net1338 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[306\] sky130_fd_sc_hd__dfrtp_1
X_16923_ _02504_ _02643_ net559 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_264_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12046_ _05928_ _05930_ _05931_ _05932_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__or4_2
XANTENNA__17218__A3 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15616__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12160__A1 game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12160__B2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19642_ clknet_leaf_15_clk game.writer.tracker.next_frame\[237\] net1289 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[237\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13417__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_284_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16854_ net1467 _02623_ _02624_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[240\]
+ sky130_fd_sc_hd__a21o_1
XANTENNA__19763__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19039__CLK net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15805_ _03416_ game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 _01817_ sky130_fd_sc_hd__nor2_1
X_19573_ clknet_leaf_49_clk game.writer.tracker.next_frame\[168\] net1294 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[168\] sky130_fd_sc_hd__dfrtp_1
X_16785_ net133 _02460_ net123 _02596_ net1833 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[198\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_87_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13997_ net940 net811 vssd1 vssd1 vccd1 vccd1 _07871_ sky130_fd_sc_hd__xor2_1
XFILLER_0_217_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_179_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18524_ net589 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_354_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12948_ net183 _06821_ _06803_ net180 vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__a211o_1
X_15736_ _01743_ _01745_ _01746_ _01747_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__or4_1
XANTENNA__09864__B1 game.CPU.applesa.ab.absxs.body_y\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18455_ net654 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__inv_2
X_12879_ game.writer.tracker.frame\[44\] game.writer.tracker.frame\[45\] net1002 vssd1
+ vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15667_ _01669_ _01672_ _01677_ _01678_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__or4_1
XFILLER_0_233_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17406_ game.CPU.kyle.L1.nextState\[1\] net1273 _02818_ vssd1 vssd1 vccd1 vccd1 _02836_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_346_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14618_ game.CPU.clock1.counter\[11\] game.CPU.clock1.counter\[10\] _08465_ vssd1
+ vssd1 vccd1 vccd1 _08469_ sky130_fd_sc_hd__and3_1
XFILLER_0_334_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15598_ net796 net431 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__xnor2_1
X_18386_ net619 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__inv_2
XANTENNA__15070__C game.CPU.applesa.ab.check_walls.above.walls\[98\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10495__B net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17337_ _01432_ _01579_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__and2_1
X_14549_ net1176 game.CPU.walls.abc.number_out\[2\] vssd1 vssd1 vccd1 vccd1 _08419_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17154__A2 _02693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16463__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_301_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17268_ net130 _02322_ net733 vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_299_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_287_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19196__D game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19007_ net1193 _00235_ _00678_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[52\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09919__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16219_ net189 _02229_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__nor2_1
XANTENNA__14912__A1 game.CPU.applesa.ab.XMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15079__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17199_ _02508_ net74 _02730_ net1627 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[479\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_259_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14912__B2 game.CPU.applesa.ab.XMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12055__X _05942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10529__A2 _04609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11400__A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_307_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17311__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16665__A1 _02243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_328_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08972_ game.CPU.randy.f1.state\[3\] vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__inv_2
X_19909_ clknet_leaf_21_clk game.writer.tracker.next_frame\[504\] net1318 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[504\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_282_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17209__A3 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 game.writer.control.detect4.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold29 game.CPU.applesa.normal1.number\[1\] vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09524__B game.CPU.applesa.ab.check_walls.above.walls\[121\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_279_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14428__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12231__A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16968__A2 _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10701__A2 _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17090__A1 _02322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13326__S1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout364_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13614__X _07488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09524_ net1097 game.CPU.applesa.ab.check_walls.above.walls\[121\] vssd1 vssd1 vccd1
+ vccd1 _03767_ sky130_fd_sc_hd__xor2_1
XFILLER_0_195_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_318_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12454__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18626__Q game.CPU.applesa.ab.absxs.body_y\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09455_ net1086 _03237_ game.CPU.applesa.ab.absxs.body_x\[69\] net917 vssd1 vssd1
+ vccd1 vccd1 _03698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout531_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout152_X net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09386_ net1106 game.CPU.applesa.ab.check_walls.above.walls\[160\] vssd1 vssd1 vccd1
+ vccd1 _03629_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18556__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13997__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17145__A2 _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19801__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1061_X net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10768__A2 _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1159_X net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16092__B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11717__A1 game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12914__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13001__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_197_Right_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10230_ _04416_ _04418_ _04422_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__or3b_1
XANTENNA__19951__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_238_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10161_ _03221_ game.CPU.randy.f1.state\[2\] _04344_ game.CPU.randy.f1.state\[4\]
+ game.CPU.randy.f1.state\[5\] vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__a2111o_1
Xfanout1005 net1009 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_4
Xfanout1016 net1019 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__buf_2
XFILLER_0_100_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1027 net1029 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_2
Xfanout1038 net1039 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout953_X net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10092_ _04293_ _04294_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__nand2_1
XANTENNA__14340__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1049 net1050 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_233_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13920_ net1043 game.CPU.applesa.ab.check_walls.above.walls\[155\] vssd1 vssd1 vccd1
+ vccd1 _07794_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout65_X net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14419__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13890__A1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16959__A2 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13890__B2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17081__A1 _02300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13851_ game.writer.tracker.frame\[563\] _06572_ net671 game.writer.tracker.frame\[564\]
+ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_260_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ game.writer.tracker.frame\[374\] game.writer.tracker.frame\[375\] net1012
+ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__mux2_1
XANTENNA__13524__X _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13782_ game.writer.tracker.frame\[177\] game.writer.tracker.frame\[179\] game.writer.tracker.frame\[180\]
+ game.writer.tracker.frame\[178\] net980 net1035 vssd1 vssd1 vccd1 vccd1 _07656_
+ sky130_fd_sc_hd__mux4_1
X_16570_ _02335_ net144 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__or2_2
XFILLER_0_201_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19331__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ game.CPU.applesa.ab.absxs.body_x\[46\] net319 vssd1 vssd1 vccd1 vccd1 _04884_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12733_ _06567_ _06571_ _06576_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__o21ai_4
X_15521_ net859 net699 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__nand2_1
XANTENNA__14068__A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15452_ _08903_ _01478_ _01477_ _01466_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18240_ net649 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
X_12664_ _06524_ _06525_ _06527_ _06540_ _06336_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__o311a_1
XFILLER_0_167_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14403_ game.CPU.applesa.ab.absxs.body_x\[71\] net874 net871 game.CPU.applesa.ab.absxs.body_y\[68\]
+ _08268_ vssd1 vssd1 vccd1 vccd1 _08277_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_100_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _05497_ _05498_ _05499_ _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__or4_1
XANTENNA__11405__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19481__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15383_ _08899_ _08915_ vssd1 vssd1 vccd1 vccd1 _08925_ sky130_fd_sc_hd__nand2_1
XANTENNA__13945__A2 game.CPU.applesa.ab.check_walls.above.walls\[67\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11204__B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18171_ net628 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__inv_2
XANTENNA__16283__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12595_ game.CPU.applesa.ab.absxs.body_x\[111\] net530 net524 game.CPU.applesa.ab.absxs.body_y\[109\]
+ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__a22o_1
XANTENNA__17136__A2 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17122_ net166 _02373_ net81 _02709_ net1827 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[423\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ _03267_ net1063 net951 _03331_ _08199_ vssd1 vssd1 vccd1 vccd1 _08208_ sky130_fd_sc_hd__a221o_1
X_11546_ game.CPU.applesa.ab.check_walls.above.walls\[150\] net254 vssd1 vssd1 vccd1
+ vccd1 _05435_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_269_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ _02422_ net83 _02686_ net1867 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[377\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_279_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16895__A1 _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15698__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14265_ _03301_ net963 net854 game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1
+ vccd1 vccd1 _08139_ sky130_fd_sc_hd__o22a_1
XANTENNA__16570__X _02494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_213_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11477_ net746 _05365_ _05364_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__o21ba_1
X_16004_ game.CPU.applesa.ab.absxs.body_x\[62\] net348 vssd1 vssd1 vccd1 vccd1 _02016_
+ sky130_fd_sc_hd__or2_1
X_13216_ net513 _07087_ _07089_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__a21o_1
X_10428_ game.CPU.bodymain1.main.pause_clk _04570_ _04572_ net1078 vssd1 vssd1 vccd1
+ vccd1 _04573_ sky130_fd_sc_hd__a31o_1
X_14196_ game.CPU.applesa.ab.absxs.body_x\[99\] net876 net960 _03325_ _08063_ vssd1
+ vssd1 vccd1 vccd1 _08070_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16730__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ net496 _07020_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__or2_1
XANTENNA__16647__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10359_ _04515_ _04519_ _04522_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__and3_1
XFILLER_0_209_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18003__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19944__RESET_B net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14122__A2 game.CPU.applesa.ab.check_walls.above.walls\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__B net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13078_ _06948_ _06951_ net678 vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_185_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ net642 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__inv_2
XANTENNA__13330__A0 _06704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13147__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16906_ net171 net95 vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_127_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12029_ _05538_ _05540_ _05915_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__or3_1
XANTENNA__12051__A game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_302_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17886_ net614 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__inv_2
XANTENNA__15065__C net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17072__A1 _02454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19625_ clknet_leaf_27_clk game.writer.tracker.next_frame\[220\] net1318 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[220\] sky130_fd_sc_hd__dfrtp_1
X_16837_ net131 _02377_ net142 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__and3_1
XANTENNA__12986__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16458__A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_251_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19556_ clknet_leaf_34_clk game.writer.tracker.next_frame\[151\] net1329 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[151\] sky130_fd_sc_hd__dfrtp_1
X_16768_ _02424_ net64 _02591_ net1801 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[187\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_220_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_338_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18507_ net579 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__inv_2
XANTENNA__09360__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18579__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15719_ _03241_ net272 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_200_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15081__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19487_ clknet_leaf_23_clk game.writer.tracker.next_frame\[82\] net1336 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[82\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19824__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_319_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16699_ _02298_ _02350_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_274_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_319_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_307_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09240_ game.CPU.walls.rand_wall.logic_enable vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__inv_2
X_18438_ net588 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_299_Right_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_319_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_196_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16905__B _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_346_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09171_ net814 vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__inv_2
X_18369_ net597 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17127__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14706__A _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13492__S0 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_313_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload51_A clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19974__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_315_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_302_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16886__B2 _02454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09519__B net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout112_A _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XANTENNA__14361__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap752 net753 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_287_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_285_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16640__B _02398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19204__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16638__A1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13756__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1021_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_227_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11265__A1_N game.CPU.applesa.ab.absxs.body_x\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08955_ game.CPU.apple_location2\[5\] vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__inv_2
XANTENNA__11784__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout481_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12124__A1 game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13321__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout579_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12124__B2 game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19354__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17063__A1 _02436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10686__A1 game.CPU.applesa.ab.absxs.body_y\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_270_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout746_A _04450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15272__A _00293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_357_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_296_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09507_ net1085 _03271_ _03272_ net1093 _03749_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__a221o_1
XANTENNA__09270__A game.CPU.applesa.enable_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_238_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09438_ net908 game.CPU.applesa.ab.absxs.body_y\[59\] game.CPU.applesa.ab.absxs.body_y\[56\]
+ net893 _03680_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__a221o_1
XFILLER_0_304_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_266_Right_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_352_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11024__B net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09369_ net1158 net824 vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__xor2_1
XANTENNA__17118__A2 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ net746 _05283_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__or2_1
XFILLER_0_352_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12380_ game.CPU.applesa.ab.absxs.body_y\[113\] net525 net366 game.CPU.applesa.ab.absxs.body_y\[115\]
+ _06256_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_278_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16877__A1 _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ net810 net249 vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__and2_1
XANTENNA__16877__B2 game.writer.tracker.frame\[257\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10610__B2 game.CPU.applesa.ab.absxs.body_x\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16390__X _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_327_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14050_ _07919_ _07921_ _07922_ _07923_ vssd1 vssd1 vccd1 vccd1 _07924_ sky130_fd_sc_hd__or4_1
X_11262_ _04845_ _04849_ _05150_ _05151_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__or4_1
XFILLER_0_321_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13001_ game.writer.tracker.frame\[534\] game.writer.tracker.frame\[535\] net1022
+ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_249_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16550__B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12363__A1 game.CPU.applesa.ab.absxs.body_y\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16629__B2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12363__B2 game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10213_ _04370_ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__nand2_1
XANTENNA__11975__A game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_249_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15447__A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ _05077_ _05078_ _05079_ _05082_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__or4b_1
XANTENNA__14351__A game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_262_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09445__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11694__B net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ game.CPU.randy.f1.c1.count\[6\] game.CPU.randy.f1.c1.count\[11\] _04329_
+ _04330_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__or4_1
XFILLER_0_280_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14070__B game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17740_ game.CPU.applesa.ab.count\[1\] _03099_ _03103_ vssd1 vssd1 vccd1 vccd1 _03104_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_265_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10126__B1 net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10075_ _04225_ _04270_ _04279_ _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__a211o_1
X_14952_ game.CPU.walls.rand_wall.count_luck\[7\] game.CPU.walls.rand_wall.count_luck\[5\]
+ game.CPU.walls.rand_wall.count_luck\[6\] vssd1 vssd1 vccd1 vccd1 _08729_ sky130_fd_sc_hd__or3b_1
XANTENNA__17054__A1 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10677__A1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13903_ net958 net795 vssd1 vssd1 vccd1 vccd1 _07777_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17671_ net194 _03058_ _03059_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__and3_1
X_14883_ net1134 _08428_ vssd1 vssd1 vccd1 vccd1 _08660_ sky130_fd_sc_hd__nor2_1
XFILLER_0_242_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18721__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16801__A1 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19410_ clknet_leaf_48_clk game.writer.tracker.next_frame\[5\] net1295 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15604__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_338_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16622_ net971 _02245_ net237 _02249_ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__a31o_1
X_13834_ _07706_ _07707_ net485 vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__mux2_1
XANTENNA__09180__A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19341_ clknet_leaf_69_clk game.CPU.applesa.twoapples.absxs.collision vssd1 vssd1
+ vccd1 vccd1 game.CPU.applesa.twoapples.collisions sky130_fd_sc_hd__dfxtp_1
X_13765_ game.writer.tracker.frame\[189\] net839 net674 game.writer.tracker.frame\[192\]
+ vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__o22a_1
X_16553_ _02318_ net144 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__nor2_2
XANTENNA__09295__A1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10977_ _03331_ net538 vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_202_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09295__B2 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15504_ net965 _01523_ _01526_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_186_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12716_ _06565_ _06581_ _06566_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__o21a_1
X_19272_ clknet_leaf_7_clk _00042_ _00902_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_16484_ net168 _02351_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__nand2_2
XFILLER_0_328_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16565__B1 _02490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13696_ game.writer.tracker.frame\[477\] game.writer.tracker.frame\[479\] game.writer.tracker.frame\[480\]
+ game.writer.tracker.frame\[478\] net974 net1012 vssd1 vssd1 vccd1 vccd1 _07570_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__18871__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19997__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13379__B1 _07229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_233_Right_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18223_ net665 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__inv_2
XFILLER_0_328_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15435_ _01432_ _01434_ _01440_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__or3b_2
X_12647_ _03229_ game.CPU.applesa.twoapples.absxs.next_head\[2\] net517 game.CPU.applesa.ab.absxs.body_y\[94\]
+ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14040__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17109__A2 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14040__B2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15366_ _08897_ _08907_ game.writer.updater.commands.cmd_num\[4\] _08878_ vssd1 vssd1
+ vccd1 vccd1 _08908_ sky130_fd_sc_hd__a2bb2o_1
X_18154_ net631 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12578_ _06216_ _06219_ _06220_ _06227_ _06291_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__a41o_1
XANTENNA__14245__B net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17105_ _02574_ net81 _02704_ net1846 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[411\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14317_ game.CPU.applesa.ab.absxs.body_x\[57\] net1066 vssd1 vssd1 vccd1 vccd1 _08191_
+ sky130_fd_sc_hd__or2_1
X_11529_ game.CPU.applesa.ab.check_walls.above.walls\[44\] net253 vssd1 vssd1 vccd1
+ vccd1 _05418_ sky130_fd_sc_hd__xnor2_1
X_15297_ game.CPU.applesa.twomode.number\[5\] _08842_ vssd1 vssd1 vccd1 vccd1 _08846_
+ sky130_fd_sc_hd__or2_1
X_18085_ net639 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_349_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold307 game.writer.tracker.frame\[90\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold318 game.CPU.randy.f1.c1.count\[15\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 game.writer.tracker.frame\[79\] vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ net53 _02516_ net119 _02682_ net1534 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[364\]
+ sky130_fd_sc_hd__a32o_1
X_14248_ game.CPU.applesa.ab.absxs.body_y\[20\] net869 net863 game.CPU.applesa.ab.absxs.body_y\[21\]
+ _08121_ vssd1 vssd1 vccd1 vccd1 _08122_ sky130_fd_sc_hd__a221o_1
XANTENNA__16281__A1_N net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15540__A1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14343__A2 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_257_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11885__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_299_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14179_ _08045_ _08046_ _08047_ _08052_ vssd1 vssd1 vccd1 vccd1 _08053_ sky130_fd_sc_hd__or4_2
Xfanout809 game.CPU.applesa.ab.check_walls.above.walls\[86\] vssd1 vssd1 vccd1 vccd1
+ net809 sky130_fd_sc_hd__buf_2
XANTENNA__19377__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15076__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18987_ net1198 _00213_ _00658_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[32\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_237_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17938_ net657 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__inv_2
XANTENNA__17045__A1 _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11109__B net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10668__B2 game.CPU.applesa.ab.absxs.body_x\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17869_ game.writer.updater.commands.count\[15\] _03186_ vssd1 vssd1 vccd1 vccd1
+ _03189_ sky130_fd_sc_hd__nand2_1
XANTENNA__15804__B net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19608_ clknet_leaf_18_clk game.writer.tracker.next_frame\[203\] net1310 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[203\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_198_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12409__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10948__B net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19539_ clknet_leaf_32_clk game.writer.tracker.next_frame\[134\] net1301 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[134\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_315_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11125__A game.CPU.applesa.ab.absxs.body_y\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_165_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16635__B _02479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_200_Right_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09223_ game.CPU.applesa.ab.check_walls.above.walls\[171\] vssd1 vssd1 vccd1 vccd1
+ _03472_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13909__A2 game.CPU.applesa.ab.check_walls.above.walls\[121\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout327_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1069_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09154_ game.CPU.applesa.ab.check_walls.above.walls\[45\] vssd1 vssd1 vccd1 vccd1
+ _03403_ sky130_fd_sc_hd__inv_2
XFILLER_0_350_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_334_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14155__B net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16859__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_233_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09085_ game.CPU.applesa.ab.absxs.body_y\[66\] vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout115_X net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1236_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14334__A2 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout696_A net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11795__A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_203_Left_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17284__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09987_ game.CPU.apple_location2\[4\] _04208_ _04209_ net1880 vssd1 vssd1 vccd1 vccd1
+ _01377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_243_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout863_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12403__B net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18744__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10204__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13845__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12648__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17036__A1 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_335_Right_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11019__B net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15714__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19470__Q game.writer.tracker.frame\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ game.CPU.applesa.ab.check_walls.collision_down _04798_ vssd1 vssd1 vccd1
+ vccd1 _04802_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11880_ game.CPU.applesa.ab.check_walls.above.walls\[141\] net305 _05763_ _05766_
+ _05767_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_67_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10831_ game.writer.control.detect4.Q\[1\] game.writer.control.detect4.Q\[0\] vssd1
+ vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__nand2b_2
XANTENNA__11306__Y _05195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_212_Left_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_315_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_251_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13550_ game.writer.tracker.frame\[109\] game.writer.tracker.frame\[111\] game.writer.tracker.frame\[112\]
+ game.writer.tracker.frame\[110\] net967 net995 vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__mux4_1
XANTENNA__15730__A game.CPU.applesa.ab.absxs.body_x\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10762_ game.CPU.applesa.ab.absxs.body_y\[90\] _04590_ net329 game.CPU.applesa.ab.absxs.body_y\[86\]
+ vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_326_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12501_ game.CPU.applesa.ab.absxs.body_x\[61\] net379 vssd1 vssd1 vccd1 vccd1 _06378_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13481_ net478 _07145_ net681 vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__o21a_1
XFILLER_0_353_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_333_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10874__A game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10693_ game.CPU.applesa.ab.absxs.body_y\[93\] _04601_ _04709_ game.CPU.applesa.ab.absxs.body_y\[89\]
+ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16562__A3 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15220_ game.CPU.applesa.normal1.number\[0\] _08780_ net758 vssd1 vssd1 vccd1 vccd1
+ _08786_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_331_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12432_ _06307_ _06308_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_171_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11689__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14065__B game.CPU.applesa.ab.check_walls.above.walls\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13781__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15151_ net1210 net1236 game.CPU.applesa.ab.check_walls.above.walls\[179\] vssd1
+ vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12584__B2 game.CPU.applesa.ab.absxs.body_x\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12363_ game.CPU.applesa.ab.absxs.body_y\[45\] net524 net365 game.CPU.applesa.ab.absxs.body_y\[47\]
+ _06239_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_340_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14102_ net942 net818 vssd1 vssd1 vccd1 vccd1 _07976_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11314_ net744 _05197_ _05199_ net567 vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__o22a_1
XANTENNA__15522__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_210_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15082_ net1211 net1237 net801 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_221_Left_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12294_ _06176_ _06179_ _06177_ _06178_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__or4b_2
XFILLER_0_239_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13533__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14033_ net948 net797 vssd1 vssd1 vccd1 vccd1 _07907_ sky130_fd_sc_hd__xnor2_1
X_18910_ clknet_leaf_3_clk _00008_ _00594_ vssd1 vssd1 vccd1 vccd1 game.CPU.modea.Qa\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_120_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_266_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11245_ game.CPU.applesa.ab.absxs.body_x\[7\] net544 net538 game.CPU.applesa.ab.absxs.body_y\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__a22o_1
X_19890_ clknet_leaf_27_clk game.writer.tracker.next_frame\[485\] net1309 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[485\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_238_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14081__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17275__A1 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09175__A game.CPU.applesa.ab.check_walls.above.walls\[81\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_18841_ clknet_leaf_73_clk _01232_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11176_ _03235_ net544 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__nand2_1
XANTENNA__15825__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10127_ net1263 net1462 net1751 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_182_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18772_ clknet_leaf_60_clk _01189_ _00509_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[78\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13836__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15984_ game.CPU.applesa.ab.check_walls.above.walls\[65\] net474 vssd1 vssd1 vccd1
+ vccd1 _01996_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12639__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17027__A1 _02524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17723_ _03085_ _03091_ _03092_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__nor3_1
XANTENNA__09504__A2 game.CPU.applesa.ab.check_walls.above.walls\[53\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_302_Right_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10058_ _04265_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__inv_2
X_14935_ _08657_ _08676_ _08699_ vssd1 vssd1 vccd1 vccd1 _08712_ sky130_fd_sc_hd__or3b_1
XANTENNA__15624__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17578__A2 _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17654_ _03047_ _03048_ _03037_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__and3b_1
XANTENNA__15589__A1 game.CPU.applesa.ab.check_walls.above.walls\[35\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14866_ _08653_ _08654_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[15\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__15589__B2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16605_ net200 _02480_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__or2_2
X_13817_ _07689_ _07690_ net498 vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17585_ game.CPU.kyle.L1.cnt_20ms\[13\] game.CPU.kyle.L1.cnt_20ms\[11\] vssd1 vssd1
+ vccd1 vccd1 _03006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_225_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14797_ game.CPU.randy.counter1.count\[7\] game.CPU.randy.counter1.count\[6\] _08608_
+ vssd1 vssd1 vccd1 vccd1 _08612_ sky130_fd_sc_hd__and3_1
XFILLER_0_175_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19324_ net1165 _01348_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twomode.counter_normal
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16536_ net202 net146 _02386_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_106_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_271_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13748_ game.writer.tracker.frame\[169\] game.writer.tracker.frame\[171\] game.writer.tracker.frame\[172\]
+ game.writer.tracker.frame\[170\] net966 net990 vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19255_ clknet_leaf_66_clk _01323_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.count_luck\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__18724__Q game.CPU.applesa.ab.absxs.body_x\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16467_ net197 _02376_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_193_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13447__S0 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13679_ net500 _07549_ _07550_ vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18617__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18206_ net666 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__inv_2
X_15418_ _08881_ _01436_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_135_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19186_ clknet_leaf_5_clk _01305_ _00848_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_331_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_310_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16398_ net172 _02280_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__or2_4
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13772__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18137_ net630 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__inv_2
X_15349_ game.writer.updater.commands.count\[11\] game.writer.updater.commands.count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _08891_ sky130_fd_sc_hd__or2_1
XANTENNA__09440__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10586__B1 _04594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09440__B2 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_269_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 game.CPU.applesa.apple_location2_n\[7\] vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 game.writer.tracker.frame\[331\] vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09637__X _03880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_257_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold126 game.writer.tracker.frame\[175\] vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18068_ net642 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__inv_2
Xhold137 game.writer.tracker.frame\[435\] vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_269_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold148 game.writer.tracker.frame\[147\] vssd1 vssd1 vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18767__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17019_ _02513_ net86 _02676_ net2003 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[353\]
+ sky130_fd_sc_hd__a2bb2o_1
Xhold159 game.writer.tracker.frame\[162\] vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15087__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09910_ _04148_ _04150_ _04151_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_282_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17266__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout606 net607 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_4
X_09841_ _04078_ _04079_ _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__and3_1
Xfanout617 net618 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__buf_4
X_20030_ net1277 vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_244_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout628 net633 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__buf_4
XFILLER_0_237_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12223__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload14_A clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout639 net640 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__buf_4
XFILLER_0_336_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14141__D _08014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ net1083 _03432_ net804 net898 _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a221o_1
XANTENNA__13288__C1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17018__A1 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_321_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout277_A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13335__A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09900__C1 _04142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_206_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10510__B1 _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout444_A _08427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13686__S0 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_293_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1186_A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13460__C1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_235_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_308_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_354_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18634__Q game.CPU.applesa.ab.absxs.body_y\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout232_X net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1353_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A _06594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14004__B2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09206_ net791 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_350_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13212__C1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Left_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_301_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11302__B _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09137_ game.CPU.applesa.ab.check_walls.above.walls\[16\] vssd1 vssd1 vccd1 vccd1
+ _03386_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1141_X net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09431__A1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09431__B2 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15504__A1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14307__A2 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ game.CPU.applesa.ab.absxs.body_y\[20\] vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout980_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15709__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_288_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13069__X _06943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19692__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 game.writer.tracker.frame\[96\] vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 game.writer.tracker.frame\[72\] vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13610__S0 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17257__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_246_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11030_ game.CPU.applesa.ab.absxs.body_y\[64\] net535 vssd1 vssd1 vccd1 vccd1 _04920_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_102_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_246_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15725__A game.CPU.applesa.ab.absxs.body_x\[53\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17009__A1 _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09282__X _03527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ net219 _06631_ net276 vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09498__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09498__B2 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11317__X _05206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14720_ _08553_ _08554_ net54 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__and3b_1
XANTENNA__17940__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09442__B game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11932_ net786 net310 vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_335_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19072__CLK net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11863_ game.CPU.applesa.ab.check_walls.above.walls\[102\] net303 _05741_ _05742_
+ _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__o2111a_1
X_14651_ _04347_ _04352_ _08489_ vssd1 vssd1 vccd1 vccd1 _08490_ sky130_fd_sc_hd__nand3_1
XFILLER_0_157_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16556__A _02403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_345_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13602_ game.writer.tracker.frame\[265\] game.writer.tracker.frame\[267\] game.writer.tracker.frame\[268\]
+ game.writer.tracker.frame\[266\] net967 net996 vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__mux4_1
X_10814_ game.CPU.applesa.ab.absxs.body_y\[117\] _04702_ vssd1 vssd1 vccd1 vccd1 _04731_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_257_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__B2 game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17370_ _03196_ _02791_ _02794_ _02798_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__a22o_1
XANTENNA__13451__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14582_ game.CPU.clock1.counter\[5\] game.CPU.clock1.counter\[8\] _08443_ vssd1 vssd1
+ vccd1 vccd1 _08444_ sky130_fd_sc_hd__and3_1
X_11794_ game.CPU.applesa.ab.check_walls.above.walls\[197\] net307 net301 game.CPU.applesa.ab.check_walls.above.walls\[198\]
+ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__o22ai_1
XANTENNA__13899__B net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16275__B net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16321_ _02262_ _02313_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__nand2_1
X_13533_ game.writer.tracker.frame\[123\] net710 net673 game.writer.tracker.frame\[124\]
+ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__o22a_1
XANTENNA__10804__B2 game.CPU.applesa.ab.absxs.body_y\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10745_ net932 game.CPU.applesa.ab.absxs.body_y\[101\] net234 _04717_ vssd1 vssd1
+ vccd1 vccd1 _01040_ sky130_fd_sc_hd__a31o_1
XANTENNA__09670__A1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Left_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09670__B2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19040_ net1188 _00271_ _00711_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[85\]
+ sky130_fd_sc_hd__dfrtp_4
X_13464_ _06663_ _07098_ net705 vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_314_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16252_ net134 _02252_ net70 net718 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__o31a_1
XANTENNA__12006__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ _03287_ _04701_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_313_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15203_ net758 _08768_ _08769_ _08770_ _08771_ vssd1 vssd1 vccd1 vccd1 _08772_ sky130_fd_sc_hd__a32o_1
X_12415_ game.CPU.applesa.ab.absxs.body_y\[35\] net364 vssd1 vssd1 vccd1 vccd1 _06292_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11212__B net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13395_ net506 _07268_ _07267_ net206 vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__a211o_1
X_16183_ _02134_ _02135_ _02193_ _02194_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__or4_2
XFILLER_0_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_346_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15134_ net1209 net1235 game.CPU.applesa.ab.check_walls.above.walls\[162\] vssd1
+ vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12346_ game.CPU.applesa.ab.absxs.body_y\[39\] net368 vssd1 vssd1 vccd1 vccd1 _06223_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_140_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15619__B net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19942_ clknet_leaf_38_clk game.writer.tracker.next_frame\[537\] net1324 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[537\] sky130_fd_sc_hd__dfrtp_1
X_15065_ net1217 net1244 net806 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09617__B game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12277_ _06159_ _06160_ _06161_ _06162_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_268_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12324__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17248__A1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14016_ net1069 game.CPU.applesa.ab.check_walls.above.walls\[184\] vssd1 vssd1 vccd1
+ vccd1 _07890_ sky130_fd_sc_hd__xor2_1
X_11228_ _03251_ net412 vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__nand2_1
X_19873_ clknet_leaf_21_clk game.writer.tracker.next_frame\[468\] net1316 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[468\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_294_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_266_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Left_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11532__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18824_ clknet_leaf_1_clk _01215_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_297_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11159_ net1269 net321 vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__or2_1
XANTENNA__18011__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18755_ clknet_leaf_53_clk _01172_ _00492_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[45\]
+ sky130_fd_sc_hd__dfrtp_4
X_15967_ game.CPU.applesa.ab.absxs.body_y\[66\] net334 vssd1 vssd1 vccd1 vccd1 _01979_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__19415__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17706_ game.CPU.walls.rand_wall.count\[1\] game.CPU.walls.rand_wall.count\[0\] net1175
+ game.CPU.walls.rand_wall.count\[2\] vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_108_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16169__C _02179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_308_Left_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14918_ _08684_ _08688_ _08694_ _08691_ vssd1 vssd1 vccd1 vccd1 _08695_ sky130_fd_sc_hd__or4b_1
XANTENNA__12493__B1 game.CPU.applesa.twoapples.absxs.next_head\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_18686_ clknet_leaf_61_clk _01103_ _00423_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_357_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09894__D1 _04136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15898_ game.CPU.applesa.ab.absxs.body_x\[41\] net474 vssd1 vssd1 vccd1 vccd1 _01910_
+ sky130_fd_sc_hd__xnor2_1
X_17637_ _08800_ net194 _03038_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__and3_1
X_14849_ _08643_ _08644_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[8\]
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_331_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19565__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17568_ _04254_ _02852_ _02879_ _02987_ _02992_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_127_Left_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19307_ net1165 _00031_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.out_random_2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11599__A2 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16519_ net167 _02368_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__nor2_8
XFILLER_0_175_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17184__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17499_ _02820_ _02826_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09661__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09661__B2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19238_ clknet_leaf_17_clk _00069_ _00876_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16931__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15734__B2 game.CPU.applesa.ab.absxs.body_y\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12218__B net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_317_Left_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13745__B1 _07618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17297__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11122__B net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19169_ clknet_leaf_57_clk _01289_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count_luck\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10019__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10559__B1 _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_230_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15529__B net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10961__B net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_300_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09527__B game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12234__A game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14152__C _08024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_136_Left_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout403 game.CPU.applesa.ab.absxs.next_head\[6\] vssd1 vssd1 vccd1 vccd1 net403
+ sky130_fd_sc_hd__buf_4
XFILLER_0_111_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout414 _04811_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_4
XFILLER_0_111_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_285_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout425 _04632_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_2
XFILLER_0_347_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout394_A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 net437 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_6
X_20013_ net1277 vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XANTENNA__15545__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09824_ net1142 game.CPU.applesa.ab.absxs.body_y\[14\] vssd1 vssd1 vccd1 vccd1 _04067_
+ sky130_fd_sc_hd__xor2_1
Xfanout447 net448 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_2
Xfanout458 net459 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1101_A game.CPU.applesa.ab.snake_head_x\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout469 net470 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_326_Left_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18629__Q game.CPU.applesa.ab.absxs.body_y\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11792__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09755_ net1132 net825 vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_253_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout561_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14473__B2 game.CPU.applesa.ab.absxs.body_y\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_241_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09686_ net904 game.CPU.applesa.ab.absxs.body_y\[102\] _03927_ _03928_ _03920_ vssd1
+ vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__a221o_1
XANTENNA__19908__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10201__B net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1091_X net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16376__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_A game.CPU.applesa.ab.check_walls.above.walls\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1189_X net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18932__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout54 net55 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_2
Xfanout65 _02560_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout76 _02690_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12882__S1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10530_ game.CPU.applesa.ab.absxs.body_x\[52\] _04609_ _04637_ game.CPU.applesa.ab.absxs.body_x\[48\]
+ vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__a22o_1
XANTENNA__11313__A game.CPU.applesa.ab.check_walls.above.walls\[64\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_335_Left_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout87 net88 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_2
XFILLER_0_107_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_330_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout98 net100 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_4
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19810__RESET_B net1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17190__A3 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17394__A_N _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12128__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13736__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11032__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_323_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10461_ net1265 _04595_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_323_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_311_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12200_ net819 net419 vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16542__C _02310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ game.writer.tracker.frame\[412\] game.writer.tracker.frame\[413\] net1035
+ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__mux2_1
XANTENNA__09718__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_clk_X clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392_ net1134 _03208_ game.CPU.apple_location\[2\] net919 _04542_ vssd1 vssd1 vccd1
+ vccd1 _04544_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout983_X net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ net831 net298 net291 game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1
+ vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14161__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ _05944_ _05945_ _05946_ _05948_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__or4_1
Xhold490 game.writer.tracker.frame\[142\] vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19438__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_257_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12711__A1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ game.CPU.applesa.ab.absxs.body_x\[52\] net415 net412 game.CPU.applesa.ab.absxs.body_x\[53\]
+ _04902_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__a221o_1
XANTENNA__11983__A game.CPU.applesa.ab.check_walls.above.walls\[180\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14997__C game.CPU.applesa.ab.check_walls.above.walls\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16870_ net157 _02425_ net99 net731 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__o31a_1
XANTENNA__10722__B1 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_341_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout970 net972 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_2
Xfanout981 net982 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_216_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09453__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15821_ game.CPU.applesa.ab.absxs.body_y\[90\] net438 net471 game.CPU.applesa.ab.absxs.body_x\[89\]
+ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__a2bb2o_1
Xfanout992 net993 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__buf_2
XANTENNA__10599__A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_271_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15661__B1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18540_ net611 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__inv_2
XFILLER_0_273_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15752_ _03378_ net272 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19588__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ net231 _06835_ _06837_ net285 vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__a31o_1
XANTENNA__09876__D1 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09340__B1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14703_ _08496_ _08503_ _08513_ _08541_ vssd1 vssd1 vccd1 vccd1 _08542_ sky130_fd_sc_hd__or4b_1
XANTENNA__11207__B net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11915_ net574 _05540_ _05537_ _05536_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__a211o_1
X_18471_ net637 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__inv_2
X_15683_ _03216_ net448 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__nand2_1
X_12895_ game.writer.tracker.frame\[26\] game.writer.tracker.frame\[27\] net1037 vssd1
+ vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__mux2_1
XANTENNA__16286__A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _02775_ _02828_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__nor2_1
X_14634_ game.CPU.clock1.counter\[16\] game.CPU.clock1.counter\[17\] _08475_ vssd1
+ vssd1 vccd1 vccd1 _08479_ sky130_fd_sc_hd__and3_1
XFILLER_0_184_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11846_ game.CPU.applesa.ab.check_walls.above.walls\[52\] net394 _05733_ vssd1 vssd1
+ vccd1 vccd1 _05734_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17353_ net1258 net1259 vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_103_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_177_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ net1175 game.CPU.walls.abc.number_out\[7\] vssd1 vssd1 vccd1 vccd1 _08430_
+ sky130_fd_sc_hd__nand2_2
X_11777_ net808 net311 vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__xnor2_1
X_16304_ _02298_ _02301_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__or2_2
XANTENNA__11223__A game.CPU.applesa.ab.absxs.body_y\[38\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_299_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13516_ net277 _07389_ net246 vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__o21a_1
X_10728_ game.CPU.applesa.ab.absxs.body_y\[31\] net330 _04714_ game.CPU.applesa.ab.absxs.body_y\[27\]
+ vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__a22o_1
X_17284_ net130 _02359_ net733 vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_190_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14496_ _08369_ vssd1 vssd1 vccd1 vccd1 _08370_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_326_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_299_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19023_ net1196 _00252_ _00694_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[68\]
+ sky130_fd_sc_hd__dfrtp_4
X_16235_ _02238_ _02241_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__nand2_4
XFILLER_0_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ _07024_ _07036_ _07037_ _07038_ net514 net705 vssd1 vssd1 vccd1 vccd1 _07321_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__12753__S net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10659_ net1078 _04695_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__nor2_2
XANTENNA__14534__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload13 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload13/X sky130_fd_sc_hd__clkbuf_4
Xclkload24 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__inv_16
XFILLER_0_301_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_298_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload35 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 clkload35/X sky130_fd_sc_hd__clkbuf_4
Xclkload46 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__10005__A2 _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09628__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ net238 _07215_ _07221_ net183 vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__a31o_1
X_16166_ _01693_ _01696_ _02176_ _02177_ _01870_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__o41a_1
Xclkload57 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__inv_12
Xclkload68 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__14253__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15117_ net1207 net1230 game.CPU.applesa.ab.check_walls.above.walls\[145\] vssd1
+ vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12329_ net1162 net846 net1271 vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_58_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09347__B game.CPU.applesa.ab.absxs.body_x\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16097_ _01847_ _01848_ _02107_ _02108_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19925_ clknet_leaf_48_clk game.writer.tracker.next_frame\[520\] net1301 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[520\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_227_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15048_ net1215 net1238 game.CPU.applesa.ab.check_walls.above.walls\[76\] vssd1 vssd1
+ vccd1 vccd1 _00270_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_114_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_282_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_267_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11505__A2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19856_ clknet_leaf_20_clk game.writer.tracker.next_frame\[451\] net1315 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[451\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_282_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_305_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18805__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16444__A2 _02395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18807_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[10\] _00544_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[10\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15084__B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19787_ clknet_leaf_24_clk game.writer.tracker.next_frame\[382\] net1346 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[382\] sky130_fd_sc_hd__dfrtp_1
X_16999_ _02485_ net89 _02671_ net1969 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[338\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12501__B net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09540_ _03779_ _03780_ _03782_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__or3_1
X_18738_ clknet_leaf_16_clk _01155_ _00475_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09471_ net1128 game.CPU.applesa.ab.absxs.body_y\[95\] vssd1 vssd1 vccd1 vccd1 _03714_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__11117__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18669_ clknet_leaf_70_clk _01086_ _00406_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[95\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_203_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_290_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10956__B net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout142_A net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_305_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_178_Right_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11441__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload7 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10972__A game.CPU.applesa.ab.absxs.body_y\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout407_A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1149_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09538__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14391__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_144_Left_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11744__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_288_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16132__A1 game.CPU.applesa.ab.absxs.body_x\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_358_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1316_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16683__A2 _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_300_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout211 net218 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_4
XFILLER_0_273_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_243_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout776_A game.CPU.applesa.ab.apple_possible\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1209 net1210 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_2
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout233 _04701_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_2
Xfanout244 net245 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_4
XANTENNA__10704__B1 _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1104_X net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout255 _05207_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_2
XFILLER_0_273_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09570__B1 game.CPU.applesa.ab.absxs.body_x\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout266 _08497_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_165_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19730__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout277 net278 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16435__A2 _02395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09807_ _04048_ _04049_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__nand2_1
Xfanout288 net289 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_2
XANTENNA_fanout943_A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout299 net301 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11308__A game.CPU.applesa.ab.check_walls.above.walls\[66\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10212__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ _03977_ _03979_ _03980_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__or3_2
XANTENNA__12457__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_153_Left_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_72_clk_X clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15722__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11027__B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09873__A1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09669_ net1101 game.CPU.applesa.ab.absxs.body_x\[37\] vssd1 vssd1 vccd1 vccd1 _03912_
+ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19880__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13082__X _06956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16738__A3 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09873__B2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ game.CPU.applesa.ab.check_walls.above.walls\[163\] net761 vssd1 vssd1 vccd1
+ vccd1 _05589_ sky130_fd_sc_hd__xnor2_2
X_12680_ _06550_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_166_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_343_Left_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_328_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_254_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _05505_ _05518_ _05519_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16834__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11562_ game.CPU.applesa.ab.check_walls.above.walls\[198\] net255 net259 net780 vssd1
+ vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12146__A2_N net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14350_ game.CPU.applesa.ab.absxs.body_x\[32\] net887 net939 _03345_ vssd1 vssd1
+ vccd1 vccd1 _08224_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17163__A3 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13301_ _06745_ _06746_ net696 vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__mux2_1
X_10513_ _04176_ _04578_ _04627_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__or3_2
XANTENNA__10786__A3 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14281_ game.CPU.applesa.ab.absxs.body_y\[86\] net947 vssd1 vssd1 vccd1 vccd1 _08155_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__11978__A game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11493_ net774 _05381_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_162_Left_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13232_ game.writer.tracker.frame\[510\] game.writer.tracker.frame\[511\] net1029
+ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__mux2_1
XANTENNA__13185__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_clk_X clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16020_ _03312_ net339 vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11697__B net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ game.CPU.bodymain1.main.score\[5\] _03196_ _04577_ vssd1 vssd1 vccd1 vccd1
+ _04579_ sky130_fd_sc_hd__or3_2
XFILLER_0_311_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11735__A2 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ game.writer.tracker.frame\[186\] game.writer.tracker.frame\[187\] net1038
+ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_343_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16123__A1 game.CPU.applesa.ab.absxs.body_x\[54\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10375_ net1081 game.CPU.apple_location2\[3\] vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18828__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12114_ _05998_ _05999_ _06000_ _05997_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_352_Left_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_265_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13094_ _06964_ _06966_ net693 vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__mux2_1
X_17971_ net662 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__inv_2
XANTENNA__10106__B game.CPU.applesa.enable_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_clk_X clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19710_ clknet_leaf_32_clk game.writer.tracker.next_frame\[305\] net1286 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[305\] sky130_fd_sc_hd__dfrtp_4
X_16922_ _02427_ _02644_ _02648_ net1766 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[284\]
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_207_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12045_ game.CPU.applesa.ab.check_walls.above.walls\[109\] net387 vssd1 vssd1 vccd1
+ vccd1 _05932_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_264_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12160__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19641_ clknet_leaf_14_clk game.writer.tracker.next_frame\[236\] net1289 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[236\] sky130_fd_sc_hd__dfrtp_1
X_16853_ net132 _02396_ net143 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_171_Left_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15804_ game.CPU.applesa.ab.check_walls.above.walls\[60\] net453 vssd1 vssd1 vccd1
+ vccd1 _01816_ sky130_fd_sc_hd__xnor2_1
X_19572_ clknet_leaf_31_clk game.writer.tracker.next_frame\[167\] net1296 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[167\] sky130_fd_sc_hd__dfrtp_1
X_16784_ _02241_ net156 vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__nor2_2
X_13996_ net960 net813 vssd1 vssd1 vccd1 vccd1 _07870_ sky130_fd_sc_hd__xor2_1
XANTENNA__16287__Y _02289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18523_ net581 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__inv_2
XANTENNA_output36_A net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15735_ _01739_ _01740_ _01742_ _01744_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_179_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_354_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ net244 _06808_ _06813_ _06818_ _06820_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__a32o_1
XANTENNA__14529__A _08028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09864__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18454_ net654 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__inv_2
XANTENNA__11671__A1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15666_ _01667_ _01668_ _01670_ _01671_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__a22o_1
X_12878_ game.writer.tracker.frame\[48\] game.writer.tracker.frame\[49\] net1007 vssd1
+ vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__mux2_2
XFILLER_0_358_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17405_ game.CPU.kyle.L1.nextState\[1\] _02834_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__nor2_1
XFILLER_0_319_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_218_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ game.CPU.clock1.counter\[9\] game.CPU.clock1.counter\[10\] _08464_ game.CPU.clock1.counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _08468_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11829_ _05553_ _05555_ _05715_ _05716_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__or4_1
X_18385_ net618 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__inv_2
XFILLER_0_233_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15597_ game.CPU.applesa.ab.check_walls.above.walls\[117\] net444 vssd1 vssd1 vccd1
+ vccd1 _01609_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12049__A net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17336_ net576 _01434_ _01582_ _08912_ vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14548_ net473 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.abduyd.next_wall\[1\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__12620__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18732__Q game.CPU.applesa.ab.absxs.body_x\[114\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_70_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19603__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_299_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17267_ net70 _02403_ _02747_ net1864 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[530\]
+ sky130_fd_sc_hd__a2bb2o_1
X_14479_ _03357_ net985 net864 game.CPU.applesa.ab.absxs.body_y\[9\] _08349_ vssd1
+ vssd1 vccd1 vccd1 _08353_ sky130_fd_sc_hd__o221a_1
XFILLER_0_102_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16901__A3 _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19006_ net1195 _00234_ _00677_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[51\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_302_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16218_ net222 net244 _02227_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__or3_2
XANTENNA__14373__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09358__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15079__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17198_ _02507_ net74 _02730_ net1615 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[478\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_286_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11726__A2 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16149_ _01725_ _01730_ _01890_ _02014_ _01618_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_307_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16114__B2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14125__B1 game.CPU.applesa.ab.check_walls.above.walls\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16665__A2 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19753__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_328_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ net1260 vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__inv_2
XANTENNA__15807__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19908_ clknet_leaf_21_clk game.writer.tracker.next_frame\[503\] net1318 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[503\] sky130_fd_sc_hd__dfrtp_1
Xhold19 game.CPU.reset_button1.eD1.Q1 vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_282_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19839_ clknet_leaf_37_clk game.writer.tracker.next_frame\[434\] net1351 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[434\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_235_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10303__Y _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12231__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17090__A2 _02693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_223_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_250_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_247_Right_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_250_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_357_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09523_ net1145 net795 vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__xor2_1
XANTENNA__18907__Q game.CPU.applesa.ab.absxs.body_y\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_318_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13343__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09454_ net1140 _03303_ game.CPU.applesa.ab.absxs.body_y\[69\] net899 _03696_ vssd1
+ vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1099_A game.CPU.applesa.ab.snake_head_x\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19133__CLK net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09385_ net1106 game.CPU.applesa.ab.check_walls.above.walls\[160\] vssd1 vssd1 vccd1
+ vccd1 _03628_ sky130_fd_sc_hd__nand2_1
XANTENNA__09607__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16654__A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout145_X net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19402__RESET_B net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09607__B2 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout524_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1266_A game.CPU.applesa.ab.absxs.body_x\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_148_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11414__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11414__B2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12611__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17145__A3 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19283__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18642__Q game.CPU.applesa.ab.absxs.body_y\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_X net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14364__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout893_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12914__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1221_X net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14902__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10160_ net1260 game.CPU.randy.f1.state\[4\] _04344_ _04353_ vssd1 vssd1 vccd1 vccd1
+ _04355_ sky130_fd_sc_hd__nor4_1
XFILLER_0_238_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15717__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1006 net1009 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1017 net1018 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__clkbuf_4
X_10091_ _04284_ _04296_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__nand2_1
Xfanout1028 net1029 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1039 net1040 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__buf_2
XANTENNA__15734__A1_N game.CPU.applesa.ab.absxs.body_y\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16388__X _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12141__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13850_ net872 game.writer.tracker.frame\[574\] game.writer.tracker.frame\[575\]
+ net708 net671 vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_260_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_214_Right_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12801_ game.writer.tracker.frame\[376\] game.writer.tracker.frame\[377\] net1033
+ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__mux2_2
X_13781_ game.writer.tracker.frame\[183\] net711 net674 game.writer.tracker.frame\[184\]
+ _07654_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__o221a_1
XANTENNA__10877__A game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10993_ game.CPU.applesa.ab.absxs.body_x\[46\] net319 vssd1 vssd1 vccd1 vccd1 _04883_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__14349__A game.CPU.applesa.ab.absxs.body_x\[35\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_201_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15520_ net944 net954 net834 _01541_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__a31o_1
X_12732_ _06604_ _06605_ net500 vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14068__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_52_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _06551_ _08922_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19626__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12663_ _06439_ _06441_ _06447_ _06539_ _06244_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__o311a_2
X_14402_ game.CPU.applesa.ab.absxs.body_x\[70\] net1056 vssd1 vssd1 vccd1 vccd1 _08276_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_100_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_309_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11614_ net802 net260 _05502_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__a21bo_1
X_18170_ net628 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__inv_2
X_15382_ _08923_ vssd1 vssd1 vccd1 vccd1 _08924_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12063__D1 _05942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11405__B2 game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12594_ game.CPU.applesa.ab.absxs.body_x\[110\] net372 game.CPU.applesa.twoapples.absxs.next_head\[3\]
+ _03257_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__a22o_1
XANTENNA__13399__S net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17121_ _02370_ _02693_ net724 vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__o21a_1
XANTENNA__19297__D net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14333_ game.CPU.applesa.ab.absxs.body_x\[74\] net1055 vssd1 vssd1 vccd1 vccd1 _08207_
+ sky130_fd_sc_hd__xor2_1
X_11545_ _05427_ _05431_ _05432_ _05433_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_67_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14084__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13158__A1 game.writer.tracker.frame\[161\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17052_ net190 _02418_ net91 _02686_ game.writer.tracker.frame\[376\] vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.next_frame\[376\] sky130_fd_sc_hd__a32o_1
XANTENNA__18650__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19776__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11476_ game.CPU.applesa.ab.check_walls.above.walls\[50\] net768 vssd1 vssd1 vccd1
+ vccd1 _05365_ sky130_fd_sc_hd__xnor2_2
X_14264_ _03235_ net1046 net863 game.CPU.applesa.ab.absxs.body_y\[77\] vssd1 vssd1
+ vccd1 vccd1 _08138_ sky130_fd_sc_hd__o22a_1
XFILLER_0_162_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13253__S1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_213_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16003_ game.CPU.applesa.ab.absxs.body_x\[62\] net348 vssd1 vssd1 vccd1 vccd1 _02015_
+ sky130_fd_sc_hd__nand2_1
X_13215_ net495 _07088_ net684 vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__a21o_1
XFILLER_0_268_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10427_ _04186_ _04571_ _04567_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__mux2_1
XANTENNA__11220__B net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ game.CPU.applesa.ab.absxs.body_x\[97\] net882 net861 game.CPU.applesa.ab.absxs.body_y\[97\]
+ _08066_ vssd1 vssd1 vccd1 vccd1 _08069_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_349_Right_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14107__B1 game.CPU.applesa.ab.check_walls.above.walls\[51\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13146_ _07016_ _07018_ net689 vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10358_ game.CPU.walls.rand_wall.counter2\[1\] game.CPU.walls.rand_wall.counter2\[0\]
+ game.CPU.walls.rand_wall.counter2\[2\] vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__a21o_1
XANTENNA__09906__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10392__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15627__B net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19006__CLK net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_295_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10392__B2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15855__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13428__A net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13077_ game.writer.tracker.frame\[230\] game.writer.tracker.frame\[231\] net998
+ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17954_ net621 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__inv_2
XFILLER_0_264_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10289_ _03214_ net1430 _04473_ _04477_ vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__o31a_1
XFILLER_0_264_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_185_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16905_ net168 _02636_ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__nor2_2
X_12028_ _05535_ _05537_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_127_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_249_Left_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17885_ net637 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_302_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12051__B net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19984__RESET_B net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17072__A2 net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19624_ clknet_leaf_27_clk game.writer.tracker.next_frame\[219\] net1321 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[219\] sky130_fd_sc_hd__dfrtp_1
X_16836_ net145 _02375_ net102 _02613_ net1689 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[232\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__10695__A2 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19156__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12986__B net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_339_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_260_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09641__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19555_ clknet_leaf_34_clk game.writer.tracker.next_frame\[150\] net1329 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[150\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11890__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16767_ _02423_ net64 _02591_ net1672 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[186\]
+ sky130_fd_sc_hd__a22o_1
X_13979_ _07848_ _07849_ _07850_ _07852_ vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__a211o_1
XANTENNA__14259__A game.CPU.applesa.ab.absxs.body_y\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10787__A game.CPU.applesa.ab.absxs.body_y\[50\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_314_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09837__B2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18506_ net586 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__inv_2
XFILLER_0_244_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15718_ _01726_ _01727_ _01728_ _01729_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__or4_2
X_19486_ clknet_leaf_26_clk game.writer.tracker.next_frame\[81\] net1312 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[81\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_66_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16698_ net205 net67 net61 _02565_ net1547 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[143\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_200_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18437_ net588 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15649_ _03421_ net270 net459 game.CPU.applesa.ab.check_walls.above.walls\[75\] _01658_
+ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__o221a_1
XANTENNA__16474__A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16583__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_196_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13397__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09170_ net815 vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18368_ net597 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_258_Left_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_313_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17127__A3 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17319_ game.writer.tracker.frame\[567\] net732 _02762_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[567\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18299_ net616 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
XFILLER_0_287_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload44_A clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12226__B net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11130__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10907__A0 net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout105_A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap753 _04355_ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16099__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_316_Right_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_285_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16638__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10383__A1 net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_227_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14441__B net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ game.CPU.apple_location2\[6\] vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_267_Left_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13321__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09525__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12124__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout474_A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19654__RESET_B net1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16810__A2 _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18637__Q game.CPU.applesa.ab.absxs.body_y\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19649__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_224_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14169__A game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09506_ net1132 game.CPU.applesa.ab.absxs.body_y\[51\] vssd1 vssd1 vccd1 vccd1 _03749_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_149_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_296_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_238_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09437_ net1149 game.CPU.applesa.ab.absxs.body_y\[57\] vssd1 vssd1 vccd1 vccd1 _03680_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_325_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_276_Left_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1171_X net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout906_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1269_X net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18673__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19799__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09368_ net1110 game.CPU.applesa.ab.check_walls.above.walls\[32\] vssd1 vssd1 vccd1
+ vccd1 _03611_ sky130_fd_sc_hd__xor2_1
XFILLER_0_352_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17118__A3 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_313_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_340_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16326__A1 game.writer.tracker.frame\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09299_ _03531_ _03532_ _03535_ _03536_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_352_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16326__B2 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13012__S net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ game.CPU.applesa.ab.check_walls.above.walls\[85\] net314 vssd1 vssd1 vccd1
+ vccd1 _05219_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14337__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16877__A2 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10610__A2 _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_320_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19029__CLK net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout896_X net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_249_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15728__A game.CPU.applesa.ab.absxs.body_x\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11261_ _04846_ _04847_ _04853_ _04854_ _04855_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a221o_1
XFILLER_0_321_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13000_ game.writer.tracker.frame\[538\] game.writer.tracker.frame\[539\] net1022
+ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__mux2_1
XANTENNA__12363__A2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10212_ net891 _04368_ _04369_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_249_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11192_ game.CPU.applesa.ab.absxs.body_x\[86\] net411 net396 game.CPU.applesa.ab.absxs.body_y\[87\]
+ _05081_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_285_Left_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14351__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ _04335_ _04336_ _04337_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__or3_2
XFILLER_0_329_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_262_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19179__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10074_ _04227_ _04275_ _04280_ _04228_ _04281_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__o221ai_1
X_14951_ _08723_ _08727_ vssd1 vssd1 vccd1 vccd1 _08728_ sky130_fd_sc_hd__and2b_1
XANTENNA__16559__A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__B1 game.CPU.applesa.ab.apple_possible\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_265_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13863__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17054__A2 _02670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ net1064 _03411_ _03412_ net1055 _07775_ vssd1 vssd1 vccd1 vccd1 _07776_ sky130_fd_sc_hd__a221o_1
X_17670_ game.CPU.kyle.L1.cnt_500hz\[13\] game.CPU.kyle.L1.cnt_500hz\[14\] _03056_
+ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__nand3_1
X_14882_ _08657_ _08658_ vssd1 vssd1 vccd1 vccd1 _08659_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_50_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19395__RESET_B net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16621_ net1814 _02526_ _02527_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[104\]
+ sky130_fd_sc_hd__a21o_1
XANTENNA__16801__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13833_ game.writer.tracker.frame\[529\] game.writer.tracker.frame\[531\] game.writer.tracker.frame\[532\]
+ game.writer.tracker.frame\[530\] net977 net1006 vssd1 vssd1 vccd1 vccd1 _07707_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_338_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09819__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09819__B2 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19340_ clknet_leaf_72_clk _01356_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.count_luck\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16552_ net170 _02318_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__nor2_1
XFILLER_0_281_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13764_ net281 _07627_ _07637_ net245 vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_294_Left_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10976_ game.CPU.applesa.ab.absxs.body_y\[74\] net402 vssd1 vssd1 vccd1 vccd1 _04866_
+ sky130_fd_sc_hd__nand2_1
X_15503_ net954 _06573_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12715_ _06583_ _06587_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19271_ clknet_leaf_6_clk _00041_ _00901_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_344_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16483_ net1735 _02426_ _02431_ _02278_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[62\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15910__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__X _04796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13695_ net491 _07566_ _07567_ _07568_ net212 vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__a311o_1
XANTENNA__16565__B2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13270__X _07144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_316_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13379__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18222_ net664 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__inv_2
XFILLER_0_343_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15434_ _01432_ _01434_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__or2_1
X_12646_ _06271_ _06272_ _06273_ _06362_ _06522_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__o311a_1
XFILLER_0_304_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18153_ net631 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__inv_2
X_15365_ _08878_ _08906_ vssd1 vssd1 vccd1 vccd1 _08907_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12577_ game.CPU.applesa.ab.absxs.body_y\[67\] net365 net524 game.CPU.applesa.ab.absxs.body_y\[65\]
+ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__a2bb2o_1
X_17104_ _02343_ net72 net735 vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__o21a_1
X_14316_ game.CPU.applesa.ab.absxs.body_x\[57\] net1066 vssd1 vssd1 vccd1 vccd1 _08190_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16868__A2 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18084_ net663 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__inv_2
X_11528_ net745 _05410_ _05412_ _05415_ _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_230_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15296_ _03525_ game.CPU.applesa.twomode.number\[0\] game.CPU.applesa.twomode.number\[1\]
+ vssd1 vssd1 vccd1 vccd1 _08845_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_349_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold308 game.writer.tracker.frame\[1\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold319 game.writer.tracker.frame\[252\] vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ _02299_ _02678_ _02682_ net1675 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[363\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14247_ game.CPU.applesa.ab.absxs.body_y\[22\] net951 vssd1 vssd1 vccd1 vccd1 _08121_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__15540__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12614__X _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11459_ net828 net256 _05347_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__a21oi_1
XANTENNA__18014__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11885__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ _08049_ _08050_ _08051_ vssd1 vssd1 vccd1 vccd1 _08052_ sky130_fd_sc_hd__or3b_1
XANTENNA__12333__Y game.CPU.applesa.twoapples.absxs.next_head\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_249_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11562__B1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13129_ game.writer.tracker.frame\[134\] game.writer.tracker.frame\[135\] net1005
+ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_239_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18986_ net1202 _00212_ _00657_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_84_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_280_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17937_ net661 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__inv_2
XANTENNA__13854__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17045__A2 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17868_ game.writer.updater.commands.count\[15\] _03186_ vssd1 vssd1 vccd1 vccd1
+ _03188_ sky130_fd_sc_hd__or2_1
XANTENNA__10668__A2 _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19607_ clknet_leaf_18_clk game.writer.tracker.next_frame\[202\] net1310 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[202\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16439__C_N _08027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16819_ net56 _02439_ net103 _02605_ net2000 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[224\]
+ sky130_fd_sc_hd__a32o_1
X_17799_ _06633_ _03134_ net556 vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_198_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19538_ clknet_leaf_32_clk game.writer.tracker.next_frame\[133\] net1296 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[133\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_191_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18696__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_315_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19941__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19469_ clknet_leaf_36_clk game.writer.tracker.next_frame\[64\] net1354 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[64\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_341_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11125__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_307_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09222_ game.CPU.applesa.ab.check_walls.above.walls\[170\] vssd1 vssd1 vccd1 vccd1
+ _03471_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10964__B net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09153_ game.CPU.applesa.ab.check_walls.above.walls\[41\] vssd1 vssd1 vccd1 vccd1
+ _03402_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout222_A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12237__A game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12593__A2 game.CPU.applesa.twoapples.absxs.next_head\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16859__A2 _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ game.CPU.applesa.ab.absxs.body_y\[72\] vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_233_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10980__A game.CPU.applesa.ab.absxs.body_x\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14452__A game.CPU.applesa.ab.absxs.body_x\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1131_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout108_X net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1229_A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19321__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09546__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout591_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_256_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout689_A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17284__A2 _02359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09986_ game.CPU.apple_location2\[5\] _04208_ _04209_ net1463 vssd1 vssd1 vccd1 vccd1
+ _01378_ sky130_fd_sc_hd__a22o_1
XFILLER_0_228_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19471__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16379__A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout856_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13355__X _07229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12700__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10830_ net1275 game.CPU.speed1.Qa\[0\] _04736_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__mux2_1
XANTENNA__11608__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_251_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15730__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10761_ game.CPU.applesa.ab.absxs.body_y\[91\] _04590_ net329 game.CPU.applesa.ab.absxs.body_y\[87\]
+ vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout909_X net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12500_ _03239_ game.CPU.applesa.twoapples.absxs.next_head\[1\] vssd1 vssd1 vccd1
+ vccd1 _06377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_325_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13480_ net501 _07135_ vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__or2_1
X_10692_ game.CPU.applesa.ab.absxs.body_y\[94\] _04601_ _04709_ game.CPU.applesa.ab.absxs.body_y\[90\]
+ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13230__A0 game.writer.tracker.frame\[512\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12431_ _03227_ game.CPU.applesa.twoapples.absxs.next_head\[2\] net360 game.CPU.applesa.ab.absxs.body_y\[100\]
+ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__o22a_1
XFILLER_0_152_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_341_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_325_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17938__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_331_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_306_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15150_ net1210 net1236 game.CPU.applesa.ab.check_walls.above.walls\[178\] vssd1
+ vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__and3_1
XANTENNA__12584__A2 game.CPU.applesa.twoapples.absxs.next_head\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12362_ game.CPU.applesa.ab.absxs.body_x\[47\] net532 vssd1 vssd1 vccd1 vccd1 _06239_
+ sky130_fd_sc_hd__xnor2_1
X_14101_ net1055 _03407_ _03408_ net1047 _07974_ vssd1 vssd1 vccd1 vccd1 _07975_ sky130_fd_sc_hd__o221a_1
X_11313_ game.CPU.applesa.ab.check_walls.above.walls\[64\] net779 vssd1 vssd1 vccd1
+ vccd1 _05202_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_210_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15081_ net1211 net1237 game.CPU.applesa.ab.check_walls.above.walls\[109\] vssd1
+ vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__and3_1
X_12293_ net829 net423 vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__nor2_1
XANTENNA__15522__A2 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14362__A game.CPU.applesa.ab.absxs.body_x\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11244_ game.CPU.applesa.ab.absxs.body_x\[108\] net324 vssd1 vssd1 vccd1 vccd1 _05134_
+ sky130_fd_sc_hd__xnor2_1
X_14032_ _07901_ _07905_ vssd1 vssd1 vccd1 vccd1 _07906_ sky130_fd_sc_hd__or2_1
XANTENNA__10347__A1 _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18569__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19814__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17275__A2 _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18840_ clknet_leaf_0_clk _01231_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_11175_ game.CPU.applesa.ab.absxs.body_x\[79\] net407 vssd1 vssd1 vccd1 vccd1 _05065_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_219_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19576__RESET_B net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16483__B1 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ game.CPU.applesa.off_bc.D net1750 net1263 vssd1 vssd1 vccd1 vccd1 _04322_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18771_ clknet_leaf_60_clk _01188_ _00508_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[77\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_262_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15905__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15983_ _03417_ net345 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_182_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ game.CPU.applesa.ab.count_luck\[3\] _03089_ vssd1 vssd1 vccd1 vccd1 _03092_
+ sky130_fd_sc_hd__nor2_1
X_10057_ _04259_ _04263_ _04264_ _04260_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__o2bb2a_1
X_14934_ _08709_ _08710_ vssd1 vssd1 vccd1 vccd1 _08711_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19964__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17653_ game.CPU.kyle.L1.cnt_500hz\[6\] game.CPU.kyle.L1.cnt_500hz\[7\] _08804_ game.CPU.kyle.L1.cnt_500hz\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__a31o_1
XANTENNA__14004__A2_N game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14865_ net1703 _08651_ vssd1 vssd1 vccd1 vccd1 _08654_ sky130_fd_sc_hd__nor2_1
XANTENNA__16786__A1 _02461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15589__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_221_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload0_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16604_ net201 _02480_ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__nor2_1
XANTENNA__11226__A game.CPU.applesa.ab.absxs.body_y\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13816_ game.writer.tracker.frame\[433\] game.writer.tracker.frame\[435\] game.writer.tracker.frame\[436\]
+ game.writer.tracker.frame\[434\] net980 net1036 vssd1 vssd1 vccd1 vccd1 _07690_
+ sky130_fd_sc_hd__mux4_1
X_17584_ game.CPU.kyle.L1.cnt_20ms\[14\] game.CPU.kyle.L1.cnt_20ms\[15\] game.CPU.kyle.L1.cnt_20ms\[16\]
+ game.CPU.kyle.L1.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__and4b_1
XFILLER_0_202_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14796_ _08610_ _08611_ vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__nor2_1
X_19323_ clknet_leaf_71_clk _01347_ _00929_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.apple_location2_n\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_16535_ net1690 _02469_ _02470_ net124 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[75\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_187_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13747_ game.writer.tracker.frame\[173\] game.writer.tracker.frame\[175\] game.writer.tracker.frame\[176\]
+ game.writer.tracker.frame\[174\] net966 net991 vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__mux4_1
XANTENNA__15640__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10959_ _03355_ net535 vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_106_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_329_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19254_ clknet_leaf_57_clk _01322_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.count_luck\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16466_ _02273_ _02419_ net559 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13678_ game.writer.tracker.frame\[490\] net841 net834 game.writer.tracker.frame\[489\]
+ vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_193_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12328__Y game.CPU.applesa.twoapples.absxs.next_head\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13447__S1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18205_ net666 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__inv_2
X_15417_ game.writer.updater.commands.count\[16\] _01443_ net833 vssd1 vssd1 vccd1
+ vccd1 _01445_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_182_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12629_ _06350_ _06351_ _06469_ _06470_ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__or4_1
XFILLER_0_72_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19185_ clknet_leaf_5_clk _01304_ _00847_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16397_ net1855 net721 _02366_ _02369_ net111 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[38\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_135_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_310_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10035__B1 _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19344__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18136_ net611 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15348_ game.writer.updater.commands.count\[6\] game.writer.updater.commands.count\[5\]
+ _08888_ _08889_ game.writer.updater.commands.count\[7\] vssd1 vssd1 vccd1 vccd1
+ _08890_ sky130_fd_sc_hd__o311a_1
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10586__A1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13587__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12980__C1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18740__Q game.CPU.applesa.ab.absxs.body_x\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_13_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold105 game.writer.tracker.frame\[294\] vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
X_18067_ net642 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__inv_2
XANTENNA__16710__A1 _02491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold116 game.writer.tracker.frame\[451\] vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ _01264_ _08828_ _08832_ vssd1 vssd1 vccd1 vccd1 _08833_ sky130_fd_sc_hd__and3b_1
Xhold127 game.writer.tracker.frame\[473\] vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold138 game.writer.tracker.frame\[457\] vssd1 vssd1 vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire180_X net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17018_ net56 _02439_ net90 _02676_ net1940 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[352\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__13524__A1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold149 game.writer.tracker.frame\[364\] vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09366__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15087__B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10338__B2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19494__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12504__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_282_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_300_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09840_ net1085 _03252_ _03320_ net1142 _04082_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__o221a_1
Xfanout607 net624 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
Xfanout618 net619 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__buf_4
XFILLER_0_272_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout629 net633 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_2
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_265_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13288__B1 _07161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09771_ net1107 _03431_ game.CPU.applesa.ab.check_walls.above.walls\[100\] net892
+ _04007_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__a221o_1
X_18969_ net1199 _00143_ _00640_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13827__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_146_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_321_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11299__C1 _05044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11838__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10959__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09900__B1 _03868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16140__A2_N net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout172_A _02254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_206_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_293_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_308_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16529__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1081_A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_235_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_307_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1179_A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09205_ game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1 vssd1 vccd1 vccd1
+ _03454_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_157_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_323_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout225_X net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout604_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17023__A_N _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13763__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12566__A2 game.CPU.applesa.twoapples.absxs.next_head\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09136_ game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1 vccd1 vccd1
+ _03385_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13497__S net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12971__C1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18711__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09067_ game.CPU.applesa.ab.absxs.body_y\[21\] vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__inv_2
XANTENNA__16701__A1 _02477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19837__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1134_X net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16701__B2 game.writer.tracker.frame\[144\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold650 game.CPU.kyle.L1.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 game.writer.tracker.frame\[201\] vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_275_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout973_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17257__A2 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_246_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18861__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19987__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15725__B net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ net1136 _04196_ _04197_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__nor3_1
XFILLER_0_228_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17009__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13526__A _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12980_ net693 _06626_ _06623_ net202 vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__o211a_1
X_11931_ _05818_ _05811_ _05810_ _05812_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__and4b_1
XFILLER_0_358_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16768__A1 _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16837__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_335_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _04343_ _04344_ _04353_ _08486_ _08488_ vssd1 vssd1 vccd1 vccd1 _08489_ sky130_fd_sc_hd__o32a_1
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11862_ _05743_ _05744_ _05748_ _05749_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_16_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13601_ net223 _07474_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_358_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11057__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10813_ net936 game.CPU.applesa.ab.absxs.body_y\[114\] _04701_ _04730_ vssd1 vssd1
+ vccd1 vccd1 _00985_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_257_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ net1275 game.CPU.speed1.Qa\[2\] vssd1 vssd1 vccd1 vccd1 _08443_ sky130_fd_sc_hd__nor2_1
X_11793_ net780 net311 vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__nor2_1
XANTENNA__14357__A game.CPU.applesa.ab.absxs.body_y\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16320_ net971 net141 _02313_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__or3b_1
XFILLER_0_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ game.writer.tracker.frame\[126\] net843 net837 game.writer.tracker.frame\[125\]
+ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__o22a_1
XFILLER_0_184_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19367__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10744_ game.CPU.applesa.ab.absxs.body_y\[105\] _04658_ vssd1 vssd1 vccd1 vccd1 _04717_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10804__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16251_ net117 net160 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__nand2_1
XANTENNA__13203__A0 _07073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12006__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_326_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13463_ net684 _07093_ _07336_ net230 vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_24_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16940__A1 _02378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10675_ net935 game.CPU.applesa.ab.absxs.body_x\[114\] net233 _04704_ vssd1 vssd1
+ vccd1 vccd1 _01097_ sky130_fd_sc_hd__a31o_1
X_15202_ game.CPU.applesa.normal1.number\[5\] _08766_ net758 vssd1 vssd1 vccd1 vccd1
+ _08771_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_313_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12414_ _06283_ _06287_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__and3_1
XANTENNA__09738__X _03981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16182_ _01732_ _01733_ _01734_ _01735_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_298_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13394_ _06864_ _06880_ net679 vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_313_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15133_ net1209 net1235 game.CPU.applesa.ab.check_walls.above.walls\[161\] vssd1
+ vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__and3_1
XANTENNA__18560__Q game.CPU.applesa.ab.absxs.body_y\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12345_ game.CPU.applesa.ab.absxs.body_x\[36\] net385 vssd1 vssd1 vccd1 vccd1 _06222_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_346_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14092__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13506__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09186__A net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19941_ clknet_leaf_38_clk game.writer.tracker.next_frame\[536\] net1330 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[536\] sky130_fd_sc_hd__dfrtp_1
X_15064_ net1218 net1245 net807 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__and3_1
X_12276_ game.CPU.applesa.ab.check_walls.above.walls\[159\] net422 vssd1 vssd1 vccd1
+ vccd1 _06162_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_268_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14015_ net959 game.CPU.applesa.ab.check_walls.above.walls\[189\] vssd1 vssd1 vccd1
+ vccd1 _07889_ sky130_fd_sc_hd__xor2_1
XANTENNA__17248__A2 _02252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11227_ game.CPU.applesa.ab.absxs.body_x\[13\] net322 vssd1 vssd1 vccd1 vccd1 _05117_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__15916__A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19872_ clknet_leaf_27_clk game.writer.tracker.next_frame\[467\] net1311 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[467\] sky130_fd_sc_hd__dfrtp_1
X_18823_ clknet_leaf_1_clk _01214_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__dfxtp_1
XANTENNA__09914__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15635__B net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158_ net1269 net321 vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_297_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10109_ _04314_ game.CPU.applesa.apple_location2_n\[6\] _04311_ vssd1 vssd1 vccd1
+ vccd1 _01346_ sky130_fd_sc_hd__mux2_1
X_11089_ game.CPU.applesa.ab.absxs.body_y\[60\] net536 vssd1 vssd1 vccd1 vccd1 _04979_
+ sky130_fd_sc_hd__or2_1
X_15966_ game.CPU.applesa.ab.absxs.body_y\[64\] net453 vssd1 vssd1 vccd1 vccd1 _01978_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12340__A _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18754_ clknet_leaf_53_clk _01171_ _00491_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[44\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_234_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14917_ _08692_ _08693_ vssd1 vssd1 vccd1 vccd1 _08694_ sky130_fd_sc_hd__or2_1
X_17705_ net1485 _03075_ _03081_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_108_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13690__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16759__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15897_ game.CPU.applesa.ab.absxs.body_x\[43\] net461 vssd1 vssd1 vccd1 vccd1 _01909_
+ sky130_fd_sc_hd__xnor2_1
X_18685_ clknet_leaf_9_clk _01102_ _00422_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09894__C1 _04132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_357_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17636_ game.CPU.kyle.L1.cnt_500hz\[0\] game.CPU.kyle.L1.cnt_500hz\[1\] vssd1 vssd1
+ vccd1 vccd1 _03038_ sky130_fd_sc_hd__or2_1
X_14848_ game.CPU.randy.f1.c1.count\[7\] game.CPU.randy.f1.c1.count\[6\] _08638_ game.CPU.randy.f1.c1.count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _08644_ sky130_fd_sc_hd__a31o_1
XFILLER_0_157_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17567_ _03361_ _02856_ _02874_ _02988_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__a2111o_1
X_14779_ game.CPU.randy.counter1.count\[17\] net265 _08595_ _08599_ vssd1 vssd1 vccd1
+ vccd1 _08600_ sky130_fd_sc_hd__o22a_1
XFILLER_0_322_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16518_ game.writer.tracker.frame\[70\] _02457_ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__and2_1
X_19306_ clknet_leaf_71_clk net1432 _00921_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.off_bc.Q2
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17184__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17498_ game.CPU.luck1.Qa\[0\] _02782_ _02818_ _02925_ _02926_ vssd1 vssd1 vccd1
+ vccd1 _02927_ sky130_fd_sc_hd__a311o_1
XFILLER_0_305_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16449_ net117 net158 _02408_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__and3_1
XANTENNA__18734__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19237_ clknet_leaf_17_clk _00068_ _00875_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16931__A1 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_332_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13745__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19168_ clknet_leaf_67_clk _01288_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count_luck\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17297__B _02370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19566__Q game.writer.tracker.frame\[161\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12953__C1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18119_ net585 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_230_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19099_ net1180 _00137_ _00770_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[144\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__16695__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18884__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12234__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17239__A2 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14152__D _08025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_257_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_245_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18202__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout415 net416 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout426 _02831_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__buf_2
X_20012_ net1276 vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
X_09823_ net1111 game.CPU.applesa.ab.absxs.body_x\[12\] vssd1 vssd1 vccd1 vccd1 _04066_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__09824__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout437 _08431_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_4
Xfanout448 _08427_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16998__A1 _02483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_240_Left_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout459 net464 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_4
XANTENNA__10731__A1 game.CPU.applesa.ab.absxs.body_y\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10731__B2 game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13356__S0 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ net1132 net825 vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__or2_1
XANTENNA__12250__A game.CPU.applesa.ab.check_walls.above.walls\[119\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14473__A2 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_241_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09685_ net1102 net1266 vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__or2_1
XANTENNA__13681__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout175_X net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout554_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16376__B _02258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13659__S1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13433__A0 _06943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18645__Q game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12249__X _06135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1084_X net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout55 _08545_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_181_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10798__B2 game.CPU.applesa.ab.absxs.body_y\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_146_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_308_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout77 net78 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__buf_2
XANTENNA__11313__B net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_330_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout88 net91 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_4
Xfanout99 net100 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_4
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1251_X net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14905__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13197__C1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12539__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10460_ _04589_ _04593_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_21_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12944__C1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_311_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09119_ net1075 vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__clkinv_4
X_10391_ net1081 _03209_ _03210_ net1096 _04541_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12130_ _06014_ _06015_ _06016_ _06013_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__a211o_1
XFILLER_0_276_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16150__A2 _02044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout976_X net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14161__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14161__B2 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ game.CPU.applesa.ab.check_walls.above.walls\[198\] net289 vssd1 vssd1 vccd1
+ vccd1 _05948_ sky130_fd_sc_hd__xnor2_1
Xhold480 game.writer.tracker.frame\[220\] vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold491 game.writer.tracker.frame\[248\] vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_257_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout88_X net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11012_ game.CPU.applesa.ab.absxs.body_x\[53\] net412 net406 _03240_ vssd1 vssd1
+ vccd1 vccd1 _04902_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13527__Y _07401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11983__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10722__A1 game.CPU.applesa.ab.absxs.body_y\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_341_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15820_ net1268 net457 net438 game.CPU.applesa.ab.absxs.body_y\[90\] vssd1 vssd1
+ vccd1 vccd1 _01832_ sky130_fd_sc_hd__a2bb2o_1
Xfanout960 net982 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11328__X _05217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout971 net972 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17951__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout982 game.CPU.applesa.y\[1\] vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__buf_6
Xfanout993 net994 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_4
XANTENNA__18607__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15661__B2 game.CPU.applesa.ab.check_walls.above.walls\[49\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15751_ game.CPU.applesa.ab.check_walls.above.walls\[3\] net463 vssd1 vssd1 vccd1
+ vccd1 _01763_ sky130_fd_sc_hd__xnor2_1
X_12963_ net497 _06836_ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16567__A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14702_ game.CPU.randy.counter1.count1\[9\] _08500_ _08504_ game.CPU.randy.counter1.count1\[8\]
+ _08540_ vssd1 vssd1 vccd1 vccd1 _08541_ sky130_fd_sc_hd__o221a_1
XFILLER_0_206_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11914_ net750 _05538_ _05801_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__o21ai_1
X_18470_ net653 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__inv_2
X_15682_ game.CPU.applesa.ab.absxs.body_y\[5\] net339 vssd1 vssd1 vccd1 vccd1 _01694_
+ sky130_fd_sc_hd__nand2_1
X_12894_ game.writer.tracker.frame\[32\] game.writer.tracker.frame\[33\] net1004 vssd1
+ vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__mux2_2
XANTENNA__14216__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17421_ _02775_ _02834_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__nor2_2
XFILLER_0_206_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14633_ game.CPU.clock1.counter\[15\] game.CPU.clock1.counter\[16\] _08474_ game.CPU.clock1.counter\[17\]
+ vssd1 vssd1 vccd1 vccd1 _08478_ sky130_fd_sc_hd__a31o_1
X_11845_ game.CPU.applesa.ab.check_walls.above.walls\[52\] net394 net303 net819 vssd1
+ vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__18757__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17352_ net1258 net1259 vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__nor2_2
XANTENNA__11504__A game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14564_ net442 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.abduyd.next_wall\[6\]
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17166__A1 _02460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11776_ _03425_ net307 vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__xnor2_1
X_16303_ net196 _02301_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__or2_1
X_13515_ _07366_ _07367_ net209 vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__mux2_1
XANTENNA__11223__B net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11998__X _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17283_ net117 _02577_ _02751_ net1831 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[542\]
+ sky130_fd_sc_hd__a22o_1
X_10727_ _04646_ _04652_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__and2_1
XFILLER_0_354_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16913__A1 _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_299_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14495_ net1278 _08368_ vssd1 vssd1 vccd1 vccd1 _08369_ sky130_fd_sc_hd__or2_2
XFILLER_0_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_190_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19022_ net1202 _00251_ _00693_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[67\]
+ sky130_fd_sc_hd__dfrtp_4
X_16234_ _02237_ _02240_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__nor2_1
X_13446_ net212 _07315_ _07319_ net283 vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__o211a_1
XANTENNA__09909__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10658_ game.CPU.applesa.ab.absxs.body_x\[32\] _04696_ _04697_ game.CPU.applesa.ab.absxs.body_x\[28\]
+ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__a22o_1
Xclkload14 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload14/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__14534__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload25 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__inv_8
XFILLER_0_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload36 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__inv_6
X_16165_ _01697_ _01700_ _01701_ _01702_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__or4_1
Xclkload47 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_298_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13377_ net222 _07249_ _07250_ net282 vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__a211o_1
XANTENNA__09628__B game.CPU.applesa.ab.absxs.body_y\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10589_ game.CPU.applesa.ab.absxs.body_x\[110\] _04665_ _04666_ game.CPU.applesa.ab.absxs.body_x\[106\]
+ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__a22o_1
Xclkload58 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12335__A net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload69 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__clkinv_8
X_15116_ net1207 net1233 game.CPU.applesa.ab.check_walls.above.walls\[144\] vssd1
+ vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__and3_1
X_12328_ net370 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.absxs.next_head\[2\]
+ sky130_fd_sc_hd__clkinv_4
XFILLER_0_279_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16096_ _01843_ _01844_ _02103_ _02104_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_58_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13586__S0 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19924_ clknet_leaf_33_clk game.writer.tracker.next_frame\[519\] net1301 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[519\] sky130_fd_sc_hd__dfrtp_1
X_15047_ net1219 net1244 game.CPU.applesa.ab.check_walls.above.walls\[75\] vssd1 vssd1
+ vccd1 vccd1 _00269_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_228_Right_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12259_ game.CPU.applesa.ab.check_walls.above.walls\[165\] net547 vssd1 vssd1 vccd1
+ vccd1 _06145_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_71_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12622__X _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_46 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_188_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19855_ clknet_leaf_20_clk game.writer.tracker.next_frame\[450\] net1315 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[450\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12341__Y game.CPU.applesa.twoapples.absxs.next_head\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_305_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18806_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[9\] _00543_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[9\] sky130_fd_sc_hd__dfrtp_1
X_19786_ clknet_leaf_24_clk game.writer.tracker.next_frame\[381\] net1346 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[381\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15084__C game.CPU.applesa.ab.check_walls.above.walls\[112\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19532__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16998_ _02483_ net90 _02671_ net2042 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[337\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_290_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_250_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18737_ clknet_leaf_13_clk _01154_ _00474_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[107\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_183_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15949_ game.CPU.applesa.ab.check_walls.above.walls\[44\] net451 vssd1 vssd1 vccd1
+ vccd1 _01961_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16477__A _02254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09331__A1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09331__B2 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09470_ net903 game.CPU.applesa.ab.absxs.body_y\[94\] game.CPU.applesa.ab.absxs.body_y\[92\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__a22o_1
X_18668_ clknet_leaf_70_clk _01085_ _00405_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[94\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_333_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16601__B1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_203_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17619_ game.CPU.kyle.L1.cnt_20ms\[12\] _03027_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__and2_1
XFILLER_0_349_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19682__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18599_ clknet_leaf_64_clk _01019_ _00336_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[80\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_82_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13105__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_290_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13966__A1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13966__B2 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17157__B2 game.writer.tracker.frame\[449\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15824__A2_N net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11133__B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16904__A1 _02477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11441__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout135_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload8 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_154_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17101__A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14444__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10972__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout302_A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_288_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16132__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16683__A3 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1211_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout201 net208 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout212 net218 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1309_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_243_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout223 net232 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09554__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout671_A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 _04657_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_273_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout245 net248 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout292_X net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11901__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 net257 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_4
Xfanout267 _08452_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_2
X_09806_ net1107 _03436_ game.CPU.applesa.ab.check_walls.above.walls\[106\] net921
+ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_165_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout278 net280 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_4
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09570__B2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout289 net292 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_213_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17490__B game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ _03975_ _03976_ _03973_ _03974_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__a211o_1
XANTENNA__11308__B net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12457__A1 net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16387__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout936_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_X net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1299_X net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09668_ net1130 game.CPU.applesa.ab.absxs.body_y\[39\] vssd1 vssd1 vccd1 vccd1 _03911_
+ sky130_fd_sc_hd__or2_1
XANTENNA__16199__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14619__B net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ net926 game.CPU.applesa.ab.absxs.body_x\[75\] game.CPU.applesa.ab.absxs.body_y\[72\]
+ net895 vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_254_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ net782 net251 net315 game.CPU.applesa.ab.check_walls.above.walls\[189\] vssd1
+ vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__17148__A1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16834__B net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11043__B net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ _05445_ _05447_ _05448_ _05449_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__or4_1
XFILLER_0_135_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13300_ net230 _07173_ net285 vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10512_ net1118 net1122 net1124 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_118_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14280_ game.CPU.applesa.ab.absxs.body_y\[84\] net868 net856 game.CPU.applesa.ab.absxs.body_y\[87\]
+ _08153_ vssd1 vssd1 vccd1 vccd1 _08154_ sky130_fd_sc_hd__a221o_1
XANTENNA__11978__B net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09729__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11492_ game.CPU.applesa.ab.check_walls.above.walls\[169\] net769 vssd1 vssd1 vccd1
+ vccd1 _05381_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13231_ game.writer.tracker.frame\[508\] game.writer.tracker.frame\[509\] net1033
+ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__mux2_1
XANTENNA__19405__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10443_ game.CPU.bodymain1.main.score\[7\] game.CPU.bodymain1.main.score\[6\] net1115
+ net1116 vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__or4_4
XFILLER_0_122_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_295_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12155__A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16850__A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12393__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ game.writer.tracker.frame\[188\] game.writer.tracker.frame\[189\] net1038
+ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_343_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16123__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ net1105 game.CPU.apple_location2\[0\] vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_276_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12113_ game.CPU.applesa.ab.check_walls.above.walls\[53\] net388 vssd1 vssd1 vccd1
+ vccd1 _06000_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11994__A game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13568__S0 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13093_ game.writer.tracker.frame\[240\] game.writer.tracker.frame\[241\] net999
+ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__mux2_2
X_17970_ net663 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_265_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19555__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12145__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16921_ _02289_ _02297_ _02643_ _02648_ net1597 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[283\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_207_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12044_ _03438_ net554 vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19640_ clknet_leaf_14_clk game.writer.tracker.next_frame\[235\] net1290 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[235\] sky130_fd_sc_hd__dfrtp_1
X_16852_ _02536_ net102 net557 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__a21oi_2
Xfanout790 game.CPU.applesa.ab.check_walls.above.walls\[148\] vssd1 vssd1 vccd1 vccd1
+ net790 sky130_fd_sc_hd__buf_2
XFILLER_0_272_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15803_ _03415_ net335 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__xnor2_1
X_16783_ _02462_ net104 net558 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a21oi_2
X_19571_ clknet_leaf_32_clk game.writer.tracker.next_frame\[166\] net1294 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[166\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15913__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11218__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13645__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13995_ net1071 game.CPU.applesa.ab.check_walls.above.walls\[72\] vssd1 vssd1 vccd1
+ vccd1 _07869_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_57_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
X_15734_ game.CPU.applesa.ab.absxs.body_y\[14\] net441 net435 game.CPU.applesa.ab.absxs.body_y\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__a2bb2o_1
X_18522_ net588 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__inv_2
XANTENNA__13740__S0 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12946_ net276 _06819_ net239 vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_354_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09864__A2 game.CPU.applesa.ab.absxs.body_y\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_319_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18453_ net654 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__inv_2
X_15665_ _01673_ _01674_ _01676_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__or3_1
X_12877_ _06749_ _06750_ net505 vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11671__A2 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_276_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11234__A game.CPU.applesa.ab.absxs.body_y\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14616_ net1482 _08465_ _08467_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[10\]
+ sky130_fd_sc_hd__a21oi_1
X_17404_ game.CPU.kyle.L1.nextState\[3\] game.CPU.kyle.L1.nextState\[2\] _02772_ vssd1
+ vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__nand3_1
X_18384_ net600 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__inv_2
X_11828_ net747 _05552_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17139__A1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_218_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15596_ _01598_ _01599_ _01606_ _01607_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12049__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17335_ net576 _02767_ _02766_ vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__o21a_1
X_14547_ _03488_ _04256_ _08417_ vssd1 vssd1 vccd1 vccd1 _08418_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11423__A2 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11759_ net784 net392 _05646_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12620__A1 game.CPU.applesa.ab.absxs.body_x\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14545__A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12620__B2 game.CPU.applesa.ab.absxs.body_y\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17266_ net176 _02319_ _02747_ net1667 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[529\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14478_ game.CPU.applesa.ab.absxs.body_y\[8\] net871 net858 game.CPU.applesa.ab.absxs.body_y\[11\]
+ _08350_ vssd1 vssd1 vccd1 vccd1 _08352_ sky130_fd_sc_hd__o221a_1
XFILLER_0_153_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16217_ _02227_ net238 net203 vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__and3b_1
XFILLER_0_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19005_ net1195 _00233_ _00676_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[50\]
+ sky130_fd_sc_hd__dfrtp_4
X_13429_ net702 _07035_ _07302_ net491 vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__o211a_1
XFILLER_0_287_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17197_ _02506_ net74 _02730_ net1733 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[477\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_259_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_302_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16148_ _01760_ _01761_ _01765_ _01766_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__or4_1
XANTENNA__17311__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14551__Y game.CPU.walls.rand_wall.abduyd.next_wall\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_307_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13595__S net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14125__A1 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14125__B2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16665__A3 _02432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16079_ _02081_ _02085_ _02089_ _02090_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__or4_1
X_08970_ net1259 vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_294_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13333__C1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_227_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19907_ clknet_leaf_21_clk game.writer.tracker.next_frame\[502\] net1318 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[502\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18922__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19838_ clknet_leaf_37_clk game.writer.tracker.next_frame\[433\] net1349 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[433\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_270_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14428__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput1 en vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_4
XANTENNA__11128__B net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13636__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19769_ clknet_leaf_28_clk game.writer.tracker.next_frame\[364\] net1287 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[364\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_48_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_211_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09522_ net1082 game.CPU.applesa.ab.check_walls.above.walls\[123\] vssd1 vssd1 vccd1
+ vccd1 _03765_ sky130_fd_sc_hd__xor2_1
XFILLER_0_211_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17378__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_318_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14439__B net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ net1131 game.CPU.applesa.ab.absxs.body_y\[71\] vssd1 vssd1 vccd1 vccd1 _03696_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_160_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout252_A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11144__A game.CPU.applesa.ab.absxs.body_y\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09384_ net1089 _03466_ _03468_ net1145 vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__a22o_1
XANTENNA__16654__B _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13630__Y _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19428__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12611__A1 game.CPU.applesa.ab.absxs.body_y\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_163_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout517_A _06214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16889__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17550__A1 net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_333_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19442__RESET_B net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14364__A1 game.CPU.applesa.ab.absxs.body_x\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16670__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout305_X net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19578__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_X net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_329_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout886_A _03368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1214_X net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10301__A_N game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1007 net1008 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__clkbuf_2
X_10090_ _04283_ _04297_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__or2_1
Xfanout1018 net1019 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_4
Xfanout1029 net1041 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__buf_2
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__A1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__B2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_261_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11350__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14419__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12849__S net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_260_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ game.writer.tracker.frame\[372\] game.writer.tracker.frame\[373\] net1012
+ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__mux2_1
XANTENNA__13093__X _06967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13780_ game.writer.tracker.frame\[182\] net844 net838 game.writer.tracker.frame\[181\]
+ vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__o22a_1
XFILLER_0_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10992_ game.CPU.applesa.ab.absxs.body_x\[44\] net415 vssd1 vssd1 vccd1 vccd1 _04882_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10877__B game.CPU.applesa.ab.apple_possible\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14349__B net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12731_ _06601_ _06603_ net677 vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12850__A1 game.writer.tracker.frame\[273\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11054__A game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15450_ net859 net853 _08930_ net834 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__or4b_1
X_12662_ _06528_ _06531_ _06538_ _06479_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16564__B _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14401_ _03237_ net1050 net985 _03304_ _08274_ vssd1 vssd1 vccd1 vccd1 _08275_ sky130_fd_sc_hd__a221o_1
X_11613_ net802 net260 _05500_ _05501_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__o211a_1
X_15381_ _08904_ _08920_ vssd1 vssd1 vccd1 vccd1 _08923_ sky130_fd_sc_hd__nor2_1
XANTENNA__12063__C1 _05934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _03270_ game.CPU.applesa.twoapples.absxs.next_head\[3\] net361 game.CPU.applesa.ab.absxs.body_y\[56\]
+ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17120_ _02369_ net57 _02708_ net1928 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[422\]
+ sky130_fd_sc_hd__a22o_1
X_14332_ _08204_ _08205_ vssd1 vssd1 vccd1 vccd1 _08206_ sky130_fd_sc_hd__nand2_1
X_11544_ net742 _05429_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14084__B game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17051_ _02544_ net90 _02686_ game.writer.tracker.frame\[375\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[375\] sky130_fd_sc_hd__a22o_1
XFILLER_0_123_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_269_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15552__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14263_ game.CPU.applesa.ab.absxs.body_x\[77\] net884 net878 game.CPU.applesa.ab.absxs.body_x\[78\]
+ _08136_ vssd1 vssd1 vccd1 vccd1 _08137_ sky130_fd_sc_hd__o221a_1
XFILLER_0_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_279_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11475_ game.CPU.applesa.ab.check_walls.above.walls\[51\] net763 vssd1 vssd1 vccd1
+ vccd1 _05364_ sky130_fd_sc_hd__xor2_2
XANTENNA__16580__A _02340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_213_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16002_ _02008_ _02013_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__or2_1
X_13214_ game.writer.tracker.frame\[420\] game.writer.tracker.frame\[421\] net1024
+ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10426_ game.CPU.bodymain1.Direction\[0\] _04568_ net1261 vssd1 vssd1 vccd1 vccd1
+ _04571_ sky130_fd_sc_hd__or3b_1
XANTENNA__15908__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14194_ game.CPU.applesa.ab.absxs.body_x\[98\] net1054 vssd1 vssd1 vccd1 vccd1 _08068_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_249_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14107__A1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ _07015_ _07017_ net684 vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__mux2_1
XANTENNA__14107__B2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10357_ _04516_ _04519_ _04521_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__and3b_1
XANTENNA__12172__X _06059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13076_ game.writer.tracker.frame\[226\] game.writer.tracker.frame\[227\] net1000
+ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__mux2_1
X_17953_ net642 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__inv_2
X_10288_ net851 game.CPU.applesa.ab.good_spot_next game.CPU.applesa.ab.apple_location\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_111_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_185_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16904_ _02477_ net93 _02642_ game.writer.tracker.frame\[272\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[272\] sky130_fd_sc_hd__a22o_1
X_12027_ _03384_ net553 vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_217_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17884_ net637 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__inv_2
XFILLER_0_228_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11341__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16804__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_302_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19623_ clknet_leaf_21_clk game.writer.tracker.next_frame\[218\] net1318 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[218\] sky130_fd_sc_hd__dfrtp_1
X_16835_ net1631 _02613_ _02614_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[231\]
+ sky130_fd_sc_hd__a21o_1
XANTENNA__15643__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14099__X _07973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16280__A1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19554_ clknet_leaf_34_clk game.writer.tracker.next_frame\[149\] net1329 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[149\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13713__S0 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09641__B net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16766_ _02425_ _02561_ net737 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__o21a_1
XFILLER_0_260_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13978_ net887 game.CPU.applesa.ab.check_walls.above.walls\[80\] _03425_ net959 _07851_
+ vssd1 vssd1 vccd1 vccd1 _07852_ sky130_fd_sc_hd__a221o_1
XANTENNA__10787__B _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_338_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14259__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18505_ net601 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__inv_2
X_12929_ _06794_ _06802_ net188 vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__o21a_1
X_15717_ _03356_ net337 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__xnor2_1
X_19485_ clknet_leaf_20_clk game.writer.tracker.next_frame\[80\] net1308 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[80\] sky130_fd_sc_hd__dfrtp_1
X_16697_ _02309_ net61 _02565_ net1875 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[142\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_200_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19953__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18436_ net581 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__inv_2
X_15648_ _03421_ net270 net439 net812 _01657_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__a221o_1
XFILLER_0_346_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_196_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18367_ net597 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__inv_2
X_15579_ _03427_ net273 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_330_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_313_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10604__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17318_ net136 _02277_ _02413_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__or3_1
XANTENNA__09369__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19720__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18298_ net616 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
XANTENNA__12507__B net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11411__B net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17249_ net112 _02454_ _02743_ net1765 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[516\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_259_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14420__A1_N net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_71_clk_X clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_280_Right_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_275_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15818__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10907__A1 game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16099__A1 game.CPU.applesa.ab.absxs.body_x\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_330_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16099__B2 game.CPU.applesa.ab.absxs.body_y\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19870__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_285_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11580__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08953_ game.CPU.apple_location2\[7\] vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__inv_2
XANTENNA__16489__X _02436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09525__A1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_149_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09525__B2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1007_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12145__A2_N net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10978__A game.CPU.applesa.ab.absxs.body_x\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13704__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16810__A3 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13085__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14169__B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09505_ net1084 _03408_ _03743_ _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__a211o_1
XFILLER_0_211_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_296_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19250__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout634_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19694__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17220__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_190_Left_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_304_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_238_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09436_ net1104 game.CPU.applesa.ab.absxs.body_x\[57\] vssd1 vssd1 vccd1 vccd1 _03679_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_304_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_24_clk_X clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09367_ net1092 game.CPU.applesa.ab.check_walls.above.walls\[34\] vssd1 vssd1 vccd1
+ vccd1 _03610_ sky130_fd_sc_hd__xor2_1
XFILLER_0_240_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_50 game.writer.tracker.frame\[305\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ net1099 game.CPU.applesa.ab.check_walls.above.walls\[81\] vssd1 vssd1 vccd1
+ vccd1 _03541_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12417__B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_39_clk_X clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ _04848_ _04850_ _04851_ _04852_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__or4_1
XFILLER_0_249_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15728__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_X net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ _04380_ _04403_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__xnor2_1
X_11191_ game.CPU.applesa.ab.absxs.body_x\[85\] net414 net319 _03232_ vssd1 vssd1
+ vccd1 vccd1 _05081_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_8_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_249_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_262_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10142_ game.CPU.randy.f1.a1.count\[7\] game.CPU.randy.f1.a1.count\[5\] _04333_ _04334_
+ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__or4_1
XFILLER_0_246_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13848__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10073_ _04238_ _04274_ _04229_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__o21ai_1
X_14950_ game.CPU.walls.rand_wall.count_luck\[5\] game.CPU.walls.rand_wall.count_luck\[4\]
+ _08726_ _08724_ vssd1 vssd1 vccd1 vccd1 _08727_ sky130_fd_sc_hd__a31o_1
XANTENNA__15744__A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout70_X net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16559__B _02486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ net890 game.CPU.applesa.ab.check_walls.above.walls\[56\] _07773_ _07774_
+ _07772_ vssd1 vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__a221o_1
X_14881_ net1081 _08421_ vssd1 vssd1 vccd1 vccd1 _08658_ sky130_fd_sc_hd__and2_1
XANTENNA__10677__A3 _04701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_345_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13832_ game.writer.tracker.frame\[534\] net845 net672 game.writer.tracker.frame\[536\]
+ _07705_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__o221a_1
X_16620_ net145 net124 _02375_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__and3_1
XFILLER_0_187_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_338_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14273__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16551_ _02237_ net167 _02479_ _02480_ net726 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__o41a_2
X_13763_ net204 _07630_ _07636_ net274 vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__o211a_1
X_10975_ _03332_ net404 vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_281_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12714_ _06583_ _06587_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__xor2_1
X_15502_ _07917_ _01507_ _01523_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__or3_1
XFILLER_0_214_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16482_ net171 _02430_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__nor2_4
X_19270_ clknet_leaf_6_clk _00040_ _00900_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_13694_ net510 _07564_ _07565_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__and3_1
XANTENNA__19743__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_273_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_344_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13379__A2 _07189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15433_ _01460_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__inv_2
XFILLER_0_214_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18221_ net664 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__inv_2
X_12645_ _06394_ _06399_ _06514_ _06521_ _06512_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__o311a_2
XTAP_TAPCELL_ROW_215_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11512__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15364_ game.writer.updater.commands.cmd_num\[4\] _08905_ vssd1 vssd1 vccd1 vccd1
+ _08906_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_14_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18152_ net631 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12576_ game.CPU.applesa.ab.absxs.body_x\[7\] net531 net360 game.CPU.applesa.ab.absxs.body_y\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__a22o_1
XANTENNA__17514__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17103_ net161 _02341_ net80 _02702_ net1505 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[410\]
+ sky130_fd_sc_hd__a32o_1
X_14315_ game.CPU.applesa.ab.absxs.body_y\[58\] net953 vssd1 vssd1 vccd1 vccd1 _08189_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11231__B net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18083_ net662 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__inv_2
X_11527_ net568 _05409_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__nor2_1
XANTENNA__16868__A3 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19893__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15295_ _03525_ game.CPU.applesa.twomode.number\[0\] game.CPU.applesa.twomode.number\[1\]
+ vssd1 vssd1 vccd1 vccd1 _08844_ sky130_fd_sc_hd__or3_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12339__A0 _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_349_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17034_ _02302_ _02517_ _02634_ net713 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__o31a_1
XFILLER_0_123_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold309 game.writer.tracker.frame\[467\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_269_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09917__A net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14246_ game.CPU.applesa.ab.absxs.body_x\[20\] net1072 vssd1 vssd1 vccd1 vccd1 _08120_
+ sky130_fd_sc_hd__or2_1
XANTENNA__15638__B net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11458_ game.CPU.applesa.ab.check_walls.above.walls\[20\] net252 vssd1 vssd1 vccd1
+ vccd1 _05347_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_269_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_312_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10409_ game.CPU.randy.f1.state\[4\] game.CPU.randy.f1.state\[1\] game.CPU.randy.f1.state\[0\]
+ _04555_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__nor4_1
X_14177_ _03255_ net1077 net858 game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1
+ vccd1 vccd1 _08051_ sky130_fd_sc_hd__o22a_1
X_11389_ net783 net260 vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__or2_1
XANTENNA__19123__CLK net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13128_ game.writer.tracker.frame\[132\] game.writer.tracker.frame\[133\] net1005
+ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__mux2_1
X_18985_ net1201 _00211_ _00656_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_239_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09507__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09507__B2 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13059_ game.writer.tracker.frame\[222\] game.writer.tracker.frame\[223\] net1016
+ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__mux2_1
X_17936_ net660 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__inv_2
XANTENNA__12630__X _06507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_264_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18030__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11314__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11314__B2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__B1 game.CPU.applesa.twoapples.absxs.next_head\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout1360 net8 vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09652__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18738__Q game.CPU.applesa.ab.absxs.body_x\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17867_ _03183_ _03185_ _03187_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__and3_1
XANTENNA__19273__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_354_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19606_ clknet_leaf_18_clk game.writer.tracker.next_frame\[201\] net1315 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[201\] sky130_fd_sc_hd__dfrtp_1
X_16818_ _02508_ net105 _02605_ net1812 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[223\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_255_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15092__C game.CPU.applesa.ab.check_walls.above.walls\[120\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17798_ _06633_ _03134_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_198_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14264__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19537_ clknet_leaf_32_clk game.writer.tracker.next_frame\[132\] net1296 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[132\] sky130_fd_sc_hd__dfrtp_1
X_16749_ game.writer.tracker.frame\[174\] _02585_ vssd1 vssd1 vccd1 vccd1 _02586_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_76_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_315_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_347_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19468_ clknet_leaf_36_clk game.writer.tracker.next_frame\[63\] net1354 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[63\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_341_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ game.CPU.applesa.ab.check_walls.above.walls\[169\] vssd1 vssd1 vccd1 vccd1
+ _03470_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18419_ net627 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__inv_2
XFILLER_0_335_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_307_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19399_ clknet_leaf_1_clk _01399_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_8_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12578__B1 _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09152_ game.CPU.applesa.ab.check_walls.above.walls\[40\] vssd1 vssd1 vccd1 vccd1
+ _03401_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12237__B net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16859__A3 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13790__A2 game.writer.tracker.frame\[432\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15829__A game.CPU.applesa.ab.absxs.body_x\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09083_ game.CPU.applesa.ab.absxs.body_y\[73\] vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout215_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09827__A net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_303_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14452__B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10980__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_326_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09746__A1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11002__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09746__B2 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09985_ game.CPU.apple_location2\[6\] _04208_ _04209_ net1633 vssd1 vssd1 vccd1 vccd1
+ _01379_ sky130_fd_sc_hd__a22o_1
XANTENNA__13783__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19616__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17036__A3 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout751_A _04442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12700__B net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10501__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18640__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16795__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19766__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_315_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16395__A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1281_X net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760_ game.CPU.applesa.ab.absxs.body_y\[96\] net263 _04719_ game.CPU.applesa.ab.absxs.body_y\[92\]
+ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_251_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09419_ net1155 game.CPU.applesa.ab.absxs.body_y\[96\] vssd1 vssd1 vccd1 vccd1 _03662_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18790__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10691_ game.CPU.applesa.ab.absxs.body_y\[95\] _04601_ _04709_ game.CPU.applesa.ab.absxs.body_y\[91\]
+ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__a22o_1
XANTENNA__10647__S _04690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12428__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13023__S net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12569__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ net1266 net377 net371 game.CPU.applesa.ab.absxs.body_x\[102\] vssd1 vssd1
+ vccd1 vccd1 _06307_ sky130_fd_sc_hd__o22a_1
XFILLER_0_164_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11051__B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13781__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ game.CPU.applesa.ab.absxs.body_x\[46\] net372 vssd1 vssd1 vccd1 vccd1 _06238_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_11_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12862__S net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14100_ net985 game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1 vccd1
+ vccd1 _07974_ sky130_fd_sc_hd__xnor2_1
X_11312_ net778 _05200_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__xnor2_1
X_15080_ net1212 net1237 game.CPU.applesa.ab.check_walls.above.walls\[108\] vssd1
+ vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__and3_1
X_12292_ net829 net424 vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_210_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14362__B net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14031_ _07896_ _07902_ _07903_ _07904_ vssd1 vssd1 vccd1 vccd1 _07905_ sky130_fd_sc_hd__or4b_1
XANTENNA__13533__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11243_ _03259_ net322 vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11174_ _03301_ net404 vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19296__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13546__X _07420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16483__B2 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ net1263 net1412 _04321_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__a21oi_1
X_18770_ clknet_leaf_60_clk _01187_ _00507_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[76\]
+ sky130_fd_sc_hd__dfrtp_1
X_15982_ _01990_ _01991_ _01992_ _01993_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__or4_1
XFILLER_0_261_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_182_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17721_ game.CPU.applesa.ab.count_luck\[3\] _03089_ vssd1 vssd1 vccd1 vccd1 _03091_
+ sky130_fd_sc_hd__and2_1
X_10056_ game.CPU.applesa.twoapples.count_luck\[2\] game.CPU.applesa.twoapples.count_luck\[0\]
+ _04262_ game.CPU.applesa.twoapples.count_luck\[1\] vssd1 vssd1 vccd1 vccd1 _04264_
+ sky130_fd_sc_hd__or4b_1
X_14933_ _08701_ _08708_ vssd1 vssd1 vccd1 vccd1 _08710_ sky130_fd_sc_hd__and2_1
XANTENNA__11507__A game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17652_ game.CPU.kyle.L1.cnt_500hz\[7\] game.CPU.kyle.L1.cnt_500hz\[8\] _03044_ vssd1
+ vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__and3_1
X_14864_ game.CPU.randy.f1.c1.count\[15\] _08651_ vssd1 vssd1 vccd1 vccd1 _08653_
+ sky130_fd_sc_hd__and2_1
XANTENNA__16786__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_221_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16576__Y _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16603_ net113 net156 _02365_ net714 vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__o31a_1
XFILLER_0_225_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13815_ game.writer.tracker.frame\[437\] game.writer.tracker.frame\[439\] game.writer.tracker.frame\[440\]
+ game.writer.tracker.frame\[438\] net980 net1039 vssd1 vssd1 vccd1 vccd1 _07689_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11226__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15921__B net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14795_ game.CPU.randy.counter1.count\[6\] _08608_ net138 vssd1 vssd1 vccd1 vccd1
+ _08611_ sky130_fd_sc_hd__o21ai_1
X_17583_ game.CPU.kyle.L1.cnt_20ms\[6\] _03003_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_159_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19322_ clknet_leaf_3_clk _01346_ _00928_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.apple_location2_n\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_13746_ net186 _07582_ _07619_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__or3_1
X_16534_ net145 _02300_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__and2_1
X_10958_ game.CPU.applesa.ab.absxs.body_y\[118\] net539 vssd1 vssd1 vccd1 vccd1 _04848_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_63_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19389__Q game.CPU.applesa.ab.snake_head_x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_317_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19253_ clknet_leaf_66_clk _01321_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.count_luck\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16465_ net172 _02335_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__nor2_4
X_13677_ game.writer.tracker.frame\[491\] net709 net672 game.writer.tracker.frame\[492\]
+ vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__o22a_1
X_10889_ _04778_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__nor2_1
XANTENNA__12338__A game.CPU.applesa.ab.absxs.body_y\[38\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18204_ net664 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__inv_2
X_15416_ game.writer.updater.commands.count\[16\] _01443_ vssd1 vssd1 vccd1 vccd1
+ _01444_ sky130_fd_sc_hd__nor2_1
X_12628_ _03337_ game.CPU.applesa.twoapples.absxs.next_head\[7\] game.CPU.applesa.twoapples.absxs.next_head\[4\]
+ _03340_ _06504_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__a221o_1
XFILLER_0_344_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16396_ net172 _02368_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__nor2_8
XFILLER_0_5_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19184_ clknet_leaf_5_clk _01303_ _00846_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_182_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_310_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10035__A1 game.CPU.applesa.ab.XMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15347_ game.writer.updater.commands.count\[9\] game.writer.updater.commands.count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _08889_ sky130_fd_sc_hd__and2_1
XANTENNA__10035__B2 game.CPU.applesa.ab.XMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18135_ net611 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__inv_2
XANTENNA__09976__A1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13772__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ _03233_ game.CPU.applesa.twoapples.absxs.next_head\[1\] net517 game.CPU.applesa.ab.absxs.body_y\[86\]
+ _06435_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18025__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13509__C1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold106 game.writer.tracker.frame\[302\] vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15278_ _08818_ _08827_ vssd1 vssd1 vccd1 vccd1 _08832_ sky130_fd_sc_hd__nand2_1
XANTENNA__16171__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11896__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18066_ net642 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__inv_2
Xhold117 game.writer.tracker.frame\[502\] vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold128 game.writer.tracker.frame\[452\] vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ _02508_ net89 _02676_ net1870 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[351\]
+ sky130_fd_sc_hd__a22o_1
Xhold139 game.writer.tracker.frame\[466\] vssd1 vssd1 vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19639__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14229_ game.CPU.applesa.ab.absxs.body_x\[41\] net1064 vssd1 vssd1 vccd1 vccd1 _08103_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__12177__A1_N game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09366__B net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15087__C game.CPU.applesa.ab.check_walls.above.walls\[115\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_282_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout608 net610 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_4
Xfanout619 net623 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ net1137 _03434_ _04011_ _04012_ _04010_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__a221o_1
XANTENNA__13288__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18968_ net1200 _00132_ _00639_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18663__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19789__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_321_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17018__A3 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17919_ net602 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
XANTENNA__12520__B net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18899_ clknet_leaf_2_clk _00004_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_2
Xfanout1190 game.CPU.walls.rand_wall.good_spot vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11417__A game.CPU.applesa.ab.check_walls.above.walls\[112\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16777__A2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16486__Y _02434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10510__A2 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_233_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_206_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11136__B net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15831__B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout165_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_293_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13460__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16529__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10975__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_235_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10274__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_347_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10813__A3 _04701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout332_A game.CPU.walls.rand_wall.abduyd.next_wall\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1074_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09204_ game.CPU.applesa.ab.check_walls.above.walls\[139\] vssd1 vssd1 vccd1 vccd1
+ _03453_ sky130_fd_sc_hd__inv_2
XANTENNA__13212__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_350_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_332_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09135_ game.CPU.applesa.ab.check_walls.above.walls\[12\] vssd1 vssd1 vccd1 vccd1
+ _03384_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout120_X net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10991__A game.CPU.applesa.ab.absxs.body_x\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout218_X net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1241_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_288_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10577__A2 net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ game.CPU.applesa.ab.absxs.body_y\[29\] vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14182__B net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold640 game.writer.tracker.frame\[339\] vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold651 game.CPU.kyle.L1.cnt_500hz\[4\] vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 game.writer.tracker.frame\[6\] vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1127_X net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_246_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout966_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ game.CPU.bodymain1.Direction\[0\] _04190_ net1261 vssd1 vssd1 vccd1 vccd1
+ _04197_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_168_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14476__B1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout78_A net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09292__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13526__B _07399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09899_ _03957_ _03959_ _03784_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__o21a_1
X_11930_ _05813_ _05814_ _05816_ _05817_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__or4_1
XANTENNA__16768__A2 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16396__Y _02369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16837__B _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout921_X net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15741__B game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11046__B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ game.CPU.applesa.ab.check_walls.above.walls\[100\] net394 vssd1 vssd1 vccd1
+ vccd1 _05749_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_335_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12857__S net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13600_ _07472_ _07473_ net500 vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__mux2_1
X_10812_ game.CPU.applesa.ab.absxs.body_y\[118\] _04702_ vssd1 vssd1 vccd1 vccd1 _04730_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14580_ game.CPU.clock1.counter\[6\] _08441_ net1275 vssd1 vssd1 vccd1 vccd1 _08442_
+ sky130_fd_sc_hd__o21ba_1
XANTENNA__13451__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ net780 net311 vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_257_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14357__B net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13531_ game.writer.tracker.frame\[127\] net710 net673 game.writer.tracker.frame\[128\]
+ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10743_ net932 game.CPU.applesa.ab.absxs.body_y\[102\] net234 _04716_ vssd1 vssd1
+ vccd1 vccd1 _01041_ sky130_fd_sc_hd__a31o_1
XANTENNA__17193__A2 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16853__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11062__A game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16250_ net113 _02257_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__nor2_2
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13462_ net513 _07088_ _07335_ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__a21o_1
XFILLER_0_164_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10674_ _03286_ net233 vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__nor2_1
XFILLER_0_180_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16572__B net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15201_ game.CPU.applesa.normal1.number\[5\] _08766_ vssd1 vssd1 vccd1 vccd1 _08770_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_137_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12413_ _06284_ _06285_ _06289_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__nor3_1
XFILLER_0_125_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16181_ _01731_ _01736_ _01737_ _01738_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_209_Right_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_341_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13393_ net679 _06861_ _07266_ net485 vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15132_ net1209 net1235 game.CPU.applesa.ab.check_walls.above.walls\[160\] vssd1
+ vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__and3_1
XFILLER_0_279_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09467__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12344_ game.CPU.applesa.ab.absxs.body_x\[36\] net381 vssd1 vssd1 vccd1 vccd1 _06221_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_152_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16153__B1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_346_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14092__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19940_ clknet_leaf_38_clk game.writer.tracker.next_frame\[535\] net1330 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[535\] sky130_fd_sc_hd__dfrtp_1
X_15063_ net1218 net1247 game.CPU.applesa.ab.check_walls.above.walls\[91\] vssd1 vssd1
+ vccd1 vccd1 _00286_ sky130_fd_sc_hd__and3_1
XFILLER_0_287_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12275_ _03463_ net421 vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__nor2_1
XANTENNA__11517__A1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_268_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14014_ net1044 game.CPU.applesa.ab.check_walls.above.walls\[187\] vssd1 vssd1 vccd1
+ vccd1 _07888_ sky130_fd_sc_hd__xor2_1
X_11226_ game.CPU.applesa.ab.absxs.body_y\[12\] net535 vssd1 vssd1 vccd1 vccd1 _05116_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19871_ clknet_leaf_27_clk game.writer.tracker.next_frame\[466\] net1311 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[466\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17248__A3 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19931__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15916__B net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19797__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18822_ clknet_leaf_2_clk _01213_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11157_ _03272_ net320 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14467__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_297_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10108_ game.CPU.applesa.twoapples.y_final\[2\] _04312_ vssd1 vssd1 vccd1 vccd1 _04314_
+ sky130_fd_sc_hd__or2_1
X_18753_ clknet_leaf_59_clk _01170_ _00490_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[39\]
+ sky130_fd_sc_hd__dfrtp_4
X_11088_ game.CPU.applesa.ab.absxs.body_y\[60\] net536 vssd1 vssd1 vccd1 vccd1 _04978_
+ sky130_fd_sc_hd__nand2_1
X_15965_ game.CPU.applesa.ab.absxs.body_y\[67\] net434 vssd1 vssd1 vccd1 vccd1 _01977_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_262_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15932__A game.CPU.applesa.ab.check_walls.above.walls\[120\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17704_ game.CPU.walls.rand_wall.count\[1\] _03075_ _03080_ vssd1 vssd1 vccd1 vccd1
+ _03081_ sky130_fd_sc_hd__o21ai_1
X_10039_ _04218_ _04220_ _04226_ _04237_ _04246_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__a41o_1
X_14916_ _08414_ _08417_ _08419_ _08421_ game.CPU.walls.rand_wall.collisions vssd1
+ vssd1 vccd1 vccd1 _08693_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_108_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18684_ clknet_leaf_8_clk _01101_ _00421_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14219__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16759__A2 _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12493__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15896_ _03343_ net335 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13690__B2 game.writer.tracker.frame\[512\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_357_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09930__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17635_ game.CPU.kyle.L1.cnt_500hz\[0\] net194 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__and2b_1
XANTENNA__15651__B net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14847_ game.CPU.randy.f1.c1.count\[7\] game.CPU.randy.f1.c1.count\[6\] game.CPU.randy.f1.c1.count\[8\]
+ _08638_ vssd1 vssd1 vccd1 vccd1 _08643_ sky130_fd_sc_hd__and4_1
XANTENNA__14548__A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17566_ _02841_ _02990_ _02989_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12876__S0 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14778_ game.CPU.randy.counter1.count\[17\] net265 _08598_ game.CPU.randy.counter1.count\[16\]
+ vssd1 vssd1 vccd1 vccd1 _08599_ sky130_fd_sc_hd__a211o_1
XANTENNA__09646__B1 game.CPU.applesa.ab.check_walls.above.walls\[157\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19305_ clknet_leaf_71_clk net1412 _00920_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.off_bc.Q1
+ sky130_fd_sc_hd__dfrtp_1
X_16517_ net1920 _02457_ _02458_ net125 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[69\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11453__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13729_ _07601_ _07602_ net492 vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_329_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17497_ _02775_ _02873_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__nor2_1
XANTENNA__17184__A2 _02322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19236_ clknet_leaf_8_clk _00067_ _00874_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_116_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16448_ net203 _02407_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__nor2_2
XFILLER_0_344_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16931__A2 _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Left_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19461__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19167_ clknet_leaf_57_clk _01287_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count_luck\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_304_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16379_ net245 _02316_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__or2_2
XFILLER_0_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11756__A1 game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09377__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18118_ net582 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_230_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16144__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19098_ net1177 _00136_ _00769_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[143\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16695__A1 _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18049_ net661 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_347_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_257_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout405 game.CPU.applesa.ab.absxs.next_head\[5\] vssd1 vssd1 vccd1 vccd1 net405
+ sky130_fd_sc_hd__buf_6
Xfanout416 _04810_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__clkbuf_8
X_09822_ net1093 game.CPU.applesa.ab.absxs.body_x\[14\] vssd1 vssd1 vccd1 vccd1 _04065_
+ sky130_fd_sc_hd__xor2_1
Xfanout427 _02831_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_2
X_20011_ net1278 vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12090__X _05977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09824__B game.CPU.applesa.ab.absxs.body_y\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout438 net439 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_4
XFILLER_0_225_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout449 net451 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_4
XANTENNA__16998__A2 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ net1160 net826 vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__or2_1
XANTENNA__13356__S1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_241_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout282_A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12250__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15842__A game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09684_ net1102 net1266 vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_241_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14458__A game.CPU.applesa.ab.absxs.body_x\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout547_A net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1191_A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout168_X net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16376__C _02354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18559__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19804__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16673__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout335_X net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout56 _02354_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1077_X net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__A2 _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_312_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout67 _02393_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__buf_4
Xfanout78 net79 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout89 net90 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16392__B net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_312_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18661__Q game.CPU.applesa.ab.absxs.body_y\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14193__A game.CPU.applesa.ab.absxs.body_x\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13292__S0 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_311_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13301__S net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ game.writer.updater.commands.count\[16\] vssd1 vssd1 vccd1 vccd1 _03367_
+ sky130_fd_sc_hd__inv_2
XANTENNA__09287__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19954__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10390_ net897 game.CPU.apple_location\[5\] game.CPU.apple_location\[0\] net910 vssd1
+ vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_115_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11967__D _05854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16686__A1 _02460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14146__C1 _08019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09049_ game.CPU.applesa.ab.absxs.body_y\[84\] vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12060_ net780 net295 vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__xnor2_1
Xhold470 game.writer.tracker.frame\[38\] vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14161__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold481 game.writer.tracker.frame\[212\] vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_276_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout969_X net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ _04895_ _04896_ _04898_ _04899_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__a211o_1
Xhold492 game.CPU.kyle.L1.currentState\[3\] vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16989__A2 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10722__A2 _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout950 game.CPU.applesa.y\[2\] vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_341_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout961 net962 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__buf_4
XANTENNA__11263__A1_N game.CPU.applesa.ab.absxs.body_y\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout972 net973 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_337_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout983 net984 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__buf_4
XFILLER_0_273_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout994 net1042 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_189_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12962_ _06779_ _06782_ net689 vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__mux2_1
X_15750_ game.CPU.applesa.ab.check_walls.above.walls\[4\] net453 vssd1 vssd1 vccd1
+ vccd1 _01762_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_231_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19334__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09876__B1 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ net750 _05538_ _05540_ net574 vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__o2bb2a_1
X_14701_ _03515_ _04351_ _08539_ vssd1 vssd1 vccd1 vccd1 _08540_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_358_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12893_ game.writer.tracker.frame\[28\] game.writer.tracker.frame\[29\] net1037 vssd1
+ vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_231_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15681_ game.CPU.applesa.ab.absxs.body_y\[4\] net454 vssd1 vssd1 vccd1 vccd1 _01693_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17420_ net1243 _02841_ _02848_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__and3_1
XFILLER_0_169_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14632_ net1980 _08475_ _08477_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[16\]
+ sky130_fd_sc_hd__a21oi_1
X_11844_ net818 net312 vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__xor2_1
XFILLER_0_157_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12227__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14621__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14563_ game.CPU.walls.rand_wall.logic_enable _08428_ _08422_ vssd1 vssd1 vccd1 vccd1
+ _08429_ sky130_fd_sc_hd__a21o_4
XANTENNA__11504__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17351_ _04638_ _02780_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__and2_1
XANTENNA__19484__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11775_ net792 net305 _05656_ _05662_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17166__A2 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _06573_ net141 _02246_ _02251_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__or4_4
XFILLER_0_222_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13514_ net226 _07363_ _07387_ net284 vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__a211o_1
X_10726_ game.CPU.applesa.ab.absxs.body_y\[36\] _04642_ _04643_ game.CPU.applesa.ab.absxs.body_y\[32\]
+ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__a22o_1
X_17282_ net176 _02258_ _02348_ _02751_ net1701 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[541\]
+ sky130_fd_sc_hd__a32o_1
X_14494_ _08362_ _08365_ _08366_ _08367_ vssd1 vssd1 vccd1 vccd1 _08368_ sky130_fd_sc_hd__and4_1
XFILLER_0_326_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_190_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18571__Q game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19021_ net1196 _00250_ _00692_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[66\]
+ sky130_fd_sc_hd__dfrtp_4
X_13445_ net488 _07318_ _07317_ net227 vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__a211o_1
X_16233_ net141 _02239_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__nor2_4
XFILLER_0_82_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10835__S _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10657_ game.CPU.applesa.ab.absxs.body_x\[33\] _04696_ _04697_ game.CPU.applesa.ab.absxs.body_x\[29\]
+ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__a22o_1
XANTENNA__16388__A_N _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload15 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__09197__A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload26 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_16
XFILLER_0_140_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13376_ net687 _06694_ _07248_ net212 vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__o211a_2
XANTENNA__16126__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload37 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__inv_6
X_16164_ _01694_ _01695_ _01698_ _01699_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a22o_1
X_10588_ game.CPU.applesa.ab.absxs.body_x\[111\] _04665_ _04666_ game.CPU.applesa.ab.absxs.body_x\[107\]
+ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload48 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__inv_6
Xclkload59 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__16677__B2 _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12327_ _04232_ _04258_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__or2_1
X_15115_ net1207 net1230 game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1
+ vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16095_ _01845_ _01846_ _02105_ _02106_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__a22o_1
XFILLER_0_267_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_192_Right_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19923_ clknet_leaf_33_clk game.writer.tracker.next_frame\[518\] net1302 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[518\] sky130_fd_sc_hd__dfrtp_1
X_15046_ net1219 net1244 game.CPU.applesa.ab.check_walls.above.walls\[74\] vssd1 vssd1
+ vccd1 vccd1 _00268_ sky130_fd_sc_hd__and3_1
X_12258_ game.CPU.applesa.ab.check_walls.above.walls\[39\] net423 vssd1 vssd1 vccd1
+ vccd1 _06144_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15646__B net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14550__B _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_188_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11209_ _03296_ net403 vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11519__X _05408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19854_ clknet_leaf_35_clk game.writer.tracker.next_frame\[449\] net1345 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[449\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_76_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12189_ net794 net417 vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__and2_1
XANTENNA__12351__A game.CPU.applesa.ab.absxs.body_y\[76\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12483__A2_N net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11910__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18805_ clknet_leaf_1_clk game.CPU.clock1.next_counter\[8\] _00542_ vssd1 vssd1 vccd1
+ vccd1 game.CPU.clock1.counter\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_305_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19785_ clknet_leaf_23_clk game.writer.tracker.next_frame\[380\] net1347 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[380\] sky130_fd_sc_hd__dfrtp_1
X_16997_ _02477_ net85 _02671_ game.writer.tracker.frame\[336\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[336\] sky130_fd_sc_hd__a22o_1
XFILLER_0_247_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_267_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18736_ clknet_leaf_13_clk _01153_ _00473_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[106\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_262_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15948_ _03403_ net336 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__xnor2_1
XANTENNA__18746__Q game.CPU.applesa.ab.absxs.body_x\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_210_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18667_ clknet_leaf_70_clk _01084_ _00404_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[93\]
+ sky130_fd_sc_hd__dfrtp_4
X_15879_ _03455_ net332 vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__nor2_1
XANTENNA__18701__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19827__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_203_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17618_ _03027_ net429 _03026_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_69_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13415__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18598_ clknet_leaf_60_clk _01018_ _00335_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[75\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_82_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_290_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17549_ net1274 net428 _02825_ _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__a31o_1
XANTENNA__13966__A2 game.CPU.applesa.ab.check_walls.above.walls\[176\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12623__C1 _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16493__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17157__A2 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19977__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18851__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload67_A clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload9 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload9/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_154_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19219_ clknet_leaf_66_clk _01313_ _00858_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_location\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17101__B _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12526__A game.CPU.applesa.ab.absxs.body_x\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout128_A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12926__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11430__A game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14391__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19207__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12960__S net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10046__A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1037_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19648__RESET_B net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout497_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13351__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 net203 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout213 net218 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_243_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout224 net232 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_4
Xfanout235 _02251_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_4
XANTENNA__19357__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout246 net247 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_4
XFILLER_0_273_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10704__A2 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17093__A1 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 _05207_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_4
X_09805_ net911 game.CPU.applesa.ab.check_walls.above.walls\[104\] game.CPU.applesa.ab.check_walls.above.walls\[105\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__o22a_1
XANTENNA_input2_A gpio_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout268 _08452_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_165_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout279 net280 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_4
XANTENNA__16668__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout664_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16840__A1 _02533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ net1128 _03345_ game.CPU.applesa.ab.absxs.body_y\[33\] net898 _03978_ vssd1
+ vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__a221o_1
XFILLER_0_213_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12457__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16387__B net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ net1130 game.CPU.applesa.ab.absxs.body_y\[39\] vssd1 vssd1 vccd1 vccd1 _03910_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1194_X net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_A net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_328_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11605__A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_328_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13406__A1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ net1148 _03332_ _03333_ net1158 _03840_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11630__A2_N net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_67_Left_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_254_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16834__C net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09569__X _03812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_294_Right_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ game.CPU.applesa.ab.check_walls.above.walls\[197\] _05213_ vssd1 vssd1 vccd1
+ vccd1 _05449_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_176_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ game.CPU.applesa.ab.absxs.body_x\[68\] _04625_ _04626_ game.CPU.applesa.ab.absxs.body_x\[64\]
+ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_351_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11491_ game.CPU.applesa.ab.check_walls.above.walls\[173\] net315 vssd1 vssd1 vccd1
+ vccd1 _05380_ sky130_fd_sc_hd__xor2_1
XANTENNA__09729__B game.CPU.applesa.ab.absxs.body_x\[35\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12917__A0 _06675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ game.writer.tracker.frame\[512\] game.writer.tracker.frame\[513\] net1001
+ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__mux2_2
XFILLER_0_17_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10442_ game.CPU.bodymain1.main.score\[7\] net1114 vssd1 vssd1 vccd1 vccd1 _04577_
+ sky130_fd_sc_hd__or2_1
XANTENNA__16108__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16850__B net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12155__B net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13161_ game.writer.tracker.frame\[192\] game.writer.tracker.frame\[193\] net1038
+ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__mux2_1
XANTENNA__15747__A _03380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12393__B2 game.CPU.applesa.ab.absxs.body_y\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12870__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10373_ net1451 net847 _04206_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_343_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_76_Left_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12112_ game.CPU.applesa.ab.check_walls.above.walls\[52\] net553 vssd1 vssd1 vccd1
+ vccd1 _05999_ sky130_fd_sc_hd__or2_1
XFILLER_0_249_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13092_ game.writer.tracker.frame\[236\] game.writer.tracker.frame\[237\] net1000
+ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__mux2_1
XANTENNA__11994__B net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_265_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14370__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16920_ _02341_ _02643_ _02648_ net1600 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[282\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17962__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ _05478_ _05482_ _05929_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_207_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17084__A1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13893__B2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16851_ net1480 _02620_ _02622_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[239\]
+ sky130_fd_sc_hd__a21o_1
XANTENNA__16578__A _02301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18724__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout780 game.CPU.applesa.ab.check_walls.above.walls\[199\] vssd1 vssd1 vccd1 vccd1
+ net780 sky130_fd_sc_hd__clkbuf_4
Xfanout791 game.CPU.applesa.ab.check_walls.above.walls\[142\] vssd1 vssd1 vccd1 vccd1
+ net791 sky130_fd_sc_hd__clkbuf_4
X_15802_ _01808_ _01810_ _01813_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__or3b_4
XANTENNA__16831__B2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19570_ clknet_leaf_32_clk game.writer.tracker.next_frame\[165\] net1294 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[165\] sky130_fd_sc_hd__dfrtp_1
X_16782_ _02458_ net107 _02595_ net1817 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[197\]
+ sky130_fd_sc_hd__a22o_1
X_13994_ net1051 game.CPU.applesa.ab.check_walls.above.walls\[75\] vssd1 vssd1 vccd1
+ vccd1 _07868_ sky130_fd_sc_hd__xor2_1
X_18521_ net580 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__inv_2
X_15733_ game.CPU.applesa.ab.absxs.body_y\[14\] net441 game.CPU.walls.rand_wall.abduyd.next_wall\[7\]
+ _03318_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__a22o_1
X_12945_ _06728_ _06733_ net219 vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_354_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Left_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18452_ net652 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15664_ game.CPU.applesa.ab.check_walls.above.walls\[51\] net461 net436 game.CPU.applesa.ab.check_walls.above.walls\[55\]
+ _01675_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__a221o_1
XFILLER_0_319_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12876_ game.writer.tracker.frame\[6\] game.writer.tracker.frame\[8\] game.writer.tracker.frame\[9\]
+ game.writer.tracker.frame\[7\] net969 net1002 vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__mux4_1
XANTENNA__18874__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_276_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17403_ game.CPU.kyle.L1.nextState\[3\] game.CPU.kyle.L1.nextState\[2\] _02772_ vssd1
+ vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__and3_1
XANTENNA__11234__B net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14615_ game.CPU.clock1.counter\[10\] _08465_ net267 vssd1 vssd1 vccd1 vccd1 _08467_
+ sky130_fd_sc_hd__o21ai_1
X_18383_ net600 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__inv_2
X_11827_ net571 _05551_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__nor2_1
XANTENNA__17139__A2 _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15595_ _03400_ net446 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_218_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11959__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17334_ _08904_ _01581_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_261_Right_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14546_ net1176 game.CPU.walls.abc.number_out\[1\] vssd1 vssd1 vccd1 vccd1 _08417_
+ sky130_fd_sc_hd__nand2_2
X_11758_ net784 net392 net301 game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1
+ vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12620__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16898__A1 _02300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10709_ _03338_ net425 vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_354_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17265_ net111 _02477_ _02747_ net1954 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[528\]
+ sky130_fd_sc_hd__a22o_1
X_14477_ _03290_ net1056 net864 game.CPU.applesa.ab.absxs.body_y\[9\] _08347_ vssd1
+ vssd1 vccd1 vccd1 _08351_ sky130_fd_sc_hd__a221o_1
X_11689_ net817 net252 vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19004_ net1194 _00231_ _00675_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[49\]
+ sky130_fd_sc_hd__dfrtp_4
X_16216_ _06607_ _02226_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__nand2_4
X_13428_ net687 _06945_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__or2_1
XANTENNA__14373__A2 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17196_ _02387_ _02493_ net71 net728 vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__o31a_1
XFILLER_0_113_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_287_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_94_Left_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13359_ _07231_ _07232_ net510 vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__mux2_1
X_16147_ game.CPU.applesa.ab.check_walls.above.walls\[110\] net439 vssd1 vssd1 vccd1
+ vccd1 _02159_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_267_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14561__A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17311__A2 _02535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10395__B1 game.CPU.applesa.ab.good_collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_307_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14125__A2 game.CPU.applesa.ab.check_walls.above.walls\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16078_ _02082_ _02083_ _02086_ _02087_ _02080_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__a221o_1
XFILLER_0_328_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_229_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19906_ clknet_leaf_21_clk game.writer.tracker.next_frame\[501\] net1318 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[501\] sky130_fd_sc_hd__dfrtp_1
X_15029_ net1228 net1256 game.CPU.applesa.ab.check_walls.above.walls\[57\] vssd1 vssd1
+ vccd1 vccd1 _00249_ sky130_fd_sc_hd__and3_1
XANTENNA__15095__C game.CPU.applesa.ab.check_walls.above.walls\[123\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17075__A1 _02460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19837_ clknet_leaf_33_clk game.writer.tracker.next_frame\[432\] net1325 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[432\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11409__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16822__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13905__A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19768_ clknet_leaf_28_clk game.writer.tracker.next_frame\[363\] net1288 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[363\] sky130_fd_sc_hd__dfrtp_1
Xinput2 gpio_in[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09390__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ net1106 game.CPU.applesa.ab.check_walls.above.walls\[120\] vssd1 vssd1 vccd1
+ vccd1 _03764_ sky130_fd_sc_hd__xor2_1
XANTENNA__11723__A1_N net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18719_ clknet_leaf_69_clk _01136_ _00456_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[89\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_250_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19699_ clknet_leaf_30_clk game.writer.tracker.next_frame\[294\] net1284 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[294\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_211_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_318_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09452_ net1140 _03303_ game.CPU.applesa.ab.absxs.body_y\[68\] net893 vssd1 vssd1
+ vccd1 vccd1 _03695_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_160_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11144__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09383_ _03618_ _03621_ _03622_ _03625_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__or4_1
XANTENNA__13495__S0 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout245_A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12611__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16889__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout412_A net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17550__A2 _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1154_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11160__A game.CPU.applesa.ab.absxs.body_y\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19829__RESET_B net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14364__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13021__C1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10047__Y _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_329_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout200_X net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09565__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14190__B net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_238_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18747__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_A net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1008 net1009 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__clkbuf_4
Xfanout1019 net1041 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09543__A2 game.CPU.applesa.ab.XMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10689__A1 game.CPU.applesa.ab.absxs.body_y\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10689__B2 game.CPU.applesa.ab.absxs.body_y\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16398__A net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout60_A _02692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_260_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09719_ net1134 game.CPU.applesa.ab.absxs.body_y\[86\] vssd1 vssd1 vccd1 vccd1 _03962_
+ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10991_ game.CPU.applesa.ab.absxs.body_x\[112\] net416 vssd1 vssd1 vccd1 vccd1 _04881_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_198_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13026__S net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12730_ _06597_ _06602_ net677 vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16845__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_328_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11054__B net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12661_ _06454_ _06535_ _06536_ _06537_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__or4_2
XFILLER_0_96_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14646__A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14052__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14052__B2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14400_ game.CPU.applesa.ab.absxs.body_x\[68\] net1074 vssd1 vssd1 vccd1 vccd1 _08274_
+ sky130_fd_sc_hd__xor2_1
X_11612_ net803 net257 vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17022__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15380_ _08920_ _08921_ vssd1 vssd1 vccd1 vccd1 _08922_ sky130_fd_sc_hd__nor2_1
X_12592_ game.CPU.applesa.ab.absxs.body_y\[57\] net525 vssd1 vssd1 vccd1 vccd1 _06469_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_343_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09464__D1 net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11543_ net566 _05426_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__xnor2_1
X_14331_ game.CPU.applesa.ab.absxs.body_y\[73\] net864 net951 _03331_ vssd1 vssd1
+ vccd1 vccd1 _08205_ sky130_fd_sc_hd__o22a_1
XFILLER_0_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12166__A game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19010__Q game.CPU.applesa.ab.check_walls.above.walls\[55\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17050_ _02419_ net83 net559 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a21oi_1
X_14262_ _03236_ net1063 net873 game.CPU.applesa.ab.absxs.body_x\[79\] vssd1 vssd1
+ vccd1 vccd1 _08136_ sky130_fd_sc_hd__o22a_1
XANTENNA__19522__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15552__A1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11474_ net818 net261 vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_269_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_351_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13213_ game.writer.tracker.frame\[424\] game.writer.tracker.frame\[425\] net1023
+ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_279_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_213_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16001_ _02009_ _02010_ _02012_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__or3b_1
XANTENNA__13563__B1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10425_ _04565_ _04566_ _04569_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__or3_1
X_14193_ game.CPU.applesa.ab.absxs.body_x\[96\] net1070 vssd1 vssd1 vccd1 vccd1 _08067_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13144_ game.writer.tracker.frame\[150\] game.writer.tracker.frame\[151\] net1023
+ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__mux2_1
XANTENNA__14107__A2 game.CPU.applesa.ab.check_walls.above.walls\[50\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10356_ game.CPU.walls.rand_wall.counter2\[2\] game.CPU.walls.rand_wall.counter2\[1\]
+ game.CPU.walls.rand_wall.counter2\[0\] game.CPU.walls.rand_wall.counter2\[3\] vssd1
+ vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__a31o_1
XANTENNA__16501__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13315__B1 _07188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19672__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15855__A2 game.CPU.walls.rand_wall.abduyd.next_wall\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13075_ game.writer.tracker.frame\[228\] game.writer.tracker.frame\[229\] net1000
+ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__mux2_1
X_17952_ net613 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__inv_2
XFILLER_0_295_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10287_ net1494 _04473_ _04476_ game.CPU.applesa.ab.start_enable vssd1 vssd1 vccd1
+ vccd1 _01317_ sky130_fd_sc_hd__a22o_1
XANTENNA__13866__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17057__A1 _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16903_ net200 net67 net92 _02642_ net1516 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[271\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_185_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12026_ net830 net388 vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15924__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17883_ net637 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__inv_2
XANTENNA__16804__A1 _02328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19622_ clknet_leaf_25_clk game.writer.tracker.next_frame\[217\] net1318 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[217\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_302_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_291_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16834_ net131 net68 net142 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__and3_1
XFILLER_0_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_330_Right_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19553_ clknet_leaf_34_clk game.writer.tracker.next_frame\[148\] net1328 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[148\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16280__A2 _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16765_ _02422_ net65 _02590_ net1974 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[185\]
+ sky130_fd_sc_hd__a22o_1
X_13977_ net1061 game.CPU.applesa.ab.check_walls.above.walls\[81\] vssd1 vssd1 vccd1
+ vccd1 _07851_ sky130_fd_sc_hd__xor2_1
X_18504_ net601 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__inv_2
X_15716_ game.CPU.applesa.ab.absxs.body_y\[10\] net441 vssd1 vssd1 vccd1 vccd1 _01728_
+ sky130_fd_sc_hd__xnor2_1
X_19484_ clknet_leaf_18_clk game.writer.tracker.next_frame\[79\] net1308 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[79\] sky130_fd_sc_hd__dfrtp_1
X_12928_ _06795_ _06800_ _06801_ net276 net238 vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__o221a_1
XFILLER_0_244_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16696_ net205 _02389_ net61 _02565_ net1670 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[141\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_200_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_346_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18435_ net588 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__inv_2
X_15647_ net812 net439 net458 game.CPU.applesa.ab.check_walls.above.walls\[75\] vssd1
+ vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__a2bb2o_1
X_12859_ _06729_ _06730_ _06731_ _06732_ net480 net677 vssd1 vssd1 vccd1 vccd1 _06733_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18028__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_346_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_196_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18366_ net596 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__inv_2
XANTENNA__12054__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15578_ net807 net454 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17317_ net176 _02416_ _02761_ net1688 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[566\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19993__RESET_B net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_313_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14529_ _08028_ _08039_ vssd1 vssd1 vccd1 vccd1 _08403_ sky130_fd_sc_hd__nor2_1
XANTENNA__09470__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18297_ net620 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
XANTENNA__09369__B net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09470__B2 net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_299_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19922__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17248_ net162 _02252_ net70 net725 vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__o31a_1
XANTENNA__15543__A1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13554__A0 game.writer.tracker.frame\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17179_ _02478_ net73 _02725_ net1922 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[464\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_259_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14291__A game.CPU.applesa.ab.absxs.body_x\[54\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09385__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16099__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17296__B2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_255_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12523__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11580__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08952_ net1153 vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__inv_2
XANTENNA__17048__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15834__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout195_A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16256__C1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10540__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10978__B net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13085__A2 _06956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout362_A net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11155__A game.CPU.applesa.ab.absxs.body_x\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09504_ net900 game.CPU.applesa.ab.check_walls.above.walls\[53\] _03745_ _03746_
+ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_296_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_338_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09435_ net1095 game.CPU.applesa.ab.absxs.body_x\[58\] vssd1 vssd1 vccd1 vccd1 _03678_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_238_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10994__A game.CPU.applesa.ab.absxs.body_x\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_304_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1271_A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_X net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11442__X _05331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09366_ net1139 net822 vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__xor2_1
XFILLER_0_304_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_40 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ net1097 game.CPU.applesa.ab.check_walls.above.walls\[81\] vssd1 vssd1 vccd1
+ vccd1 _03540_ sky130_fd_sc_hd__nand2_1
XANTENNA__16681__A _02238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_51 game.writer.tracker.frame\[305\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_X net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09994__S _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14337__A2 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout996_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19695__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13640__S0 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17287__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_249_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10210_ _04400_ _04402_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_293_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11190_ game.CPU.applesa.ab.absxs.body_x\[85\] net414 net396 game.CPU.applesa.ab.absxs.body_y\[87\]
+ _05072_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_249_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ game.CPU.randy.f1.a1.count\[13\] game.CPU.randy.f1.a1.count\[12\] game.CPU.randy.f1.a1.count\[15\]
+ game.CPU.randy.f1.a1.count\[14\] vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_262_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17039__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09582__X _03825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11049__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ _04234_ _04267_ _04235_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__o21ba_1
XANTENNA__15744__B net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout951_X net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12720__Y _06594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13900_ net942 net816 vssd1 vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__or2_1
XANTENNA__09742__B net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14880_ net1081 _08421_ vssd1 vssd1 vccd1 vccd1 _08657_ sky130_fd_sc_hd__nor2_1
X_13831_ game.writer.tracker.frame\[535\] net709 net836 game.writer.tracker.frame\[533\]
+ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__o22a_1
XANTENNA__19075__CLK net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_345_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19005__Q game.CPU.applesa.ab.check_walls.above.walls\[50\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16550_ net188 net173 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__nand2_2
XFILLER_0_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13762_ net504 _07631_ _07632_ _07635_ net224 vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__a311o_1
X_10974_ game.CPU.applesa.ab.absxs.body_x\[72\] net415 vssd1 vssd1 vccd1 vccd1 _04864_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__17211__A1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15501_ net992 net853 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__nor2_1
XFILLER_0_328_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12713_ _06580_ _06586_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10834__A1 net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16481_ net198 _02308_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__or2_2
X_13693_ game.writer.tracker.frame\[506\] net843 net839 game.writer.tracker.frame\[505\]
+ vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__o22a_1
XFILLER_0_214_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_273_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18220_ net664 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__inv_2
X_15432_ _01450_ _01459_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__or2_1
XFILLER_0_344_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12644_ _06463_ _06464_ _06515_ _06518_ _06520_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__o32a_1
XFILLER_0_343_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_215_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18151_ net630 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__inv_2
X_15363_ game.writer.updater.commands.cmd_num\[1\] game.writer.updater.commands.cmd_num\[0\]
+ game.writer.updater.commands.cmd_num\[2\] game.writer.updater.commands.cmd_num\[3\]
+ vssd1 vssd1 vccd1 vccd1 _08905_ sky130_fd_sc_hd__and4_1
XFILLER_0_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12575_ _03226_ net384 vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09452__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18912__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09452__B2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17514__A2 _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17102_ net1654 _02702_ _02703_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[409\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_230_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14314_ game.CPU.applesa.ab.absxs.body_y\[58\] net953 vssd1 vssd1 vccd1 vccd1 _08188_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18082_ net663 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__inv_2
X_11526_ net779 _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16722__B1 _02576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15919__B net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15294_ _00029_ _08840_ _08841_ _08843_ vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__o22a_1
XFILLER_0_230_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_349_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17033_ _02533_ net91 _02681_ net1486 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[362\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_351_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11457_ _05342_ _05343_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__and3_1
X_14245_ game.CPU.applesa.ab.absxs.body_x\[20\] net1072 vssd1 vssd1 vccd1 vccd1 _08119_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__09917__B _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17278__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10408_ game.CPU.randy.f1.state\[3\] game.CPU.randy.f1.state\[2\] vssd1 vssd1 vccd1
+ vccd1 _04555_ sky130_fd_sc_hd__or2_1
XFILLER_0_256_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14176_ _03255_ net1074 net883 game.CPU.applesa.ab.absxs.body_x\[105\] vssd1 vssd1
+ vccd1 vccd1 _08050_ sky130_fd_sc_hd__a22o_1
X_11388_ net783 net260 vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__nand2_1
XANTENNA__12343__B net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13127_ game.writer.tracker.frame\[136\] game.writer.tracker.frame\[137\] net1005
+ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__mux2_1
X_10339_ net1644 _04508_ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__xnor2_1
X_18984_ net1197 _00209_ _00655_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_226_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ game.writer.tracker.frame\[218\] game.writer.tracker.frame\[219\] net1016
+ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__mux2_1
X_17935_ net660 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__inv_2
XFILLER_0_280_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19418__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__A1 game.CPU.applesa.ab.absxs.body_x\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1350 net1351 vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__clkbuf_2
X_12009_ game.CPU.applesa.ab.check_walls.above.walls\[77\] net388 vssd1 vssd1 vccd1
+ vccd1 _05896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_264_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17866_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__inv_2
XANTENNA__09652__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19605_ clknet_leaf_20_clk game.writer.tracker.next_frame\[200\] net1317 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[200\] sky130_fd_sc_hd__dfrtp_1
X_16817_ _02507_ net105 _02605_ net1648 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[222\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_255_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17797_ _01532_ _03134_ _03137_ net721 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14264__B2 game.CPU.applesa.ab.absxs.body_y\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_198_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_347_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19536_ clknet_leaf_32_clk game.writer.tracker.next_frame\[131\] net1291 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[131\] sky130_fd_sc_hd__dfrtp_1
X_16748_ _02394_ net98 net718 vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__o21a_1
XANTENNA__19568__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14557__Y _08425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_315_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18754__Q game.CPU.applesa.ab.absxs.body_x\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19467_ clknet_leaf_39_clk game.writer.tracker.next_frame\[62\] net1358 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[62\] sky130_fd_sc_hd__dfrtp_1
X_16679_ net173 _02237_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__or2_1
X_09220_ game.CPU.applesa.ab.check_walls.above.walls\[168\] vssd1 vssd1 vccd1 vccd1
+ _03469_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18418_ net627 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__inv_2
XFILLER_0_185_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19398_ clknet_leaf_47_clk game.writer.control.next\[1\] net1298 vssd1 vssd1 vccd1
+ vccd1 game.writer.control.current\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12518__B net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13775__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18592__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09151_ net823 vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__inv_2
X_18349_ net594 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14319__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09082_ game.CPU.applesa.ab.absxs.body_y\[74\] vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__inv_2
XANTENNA__15829__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_342_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_287_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09827__B game.CPU.applesa.ab.absxs.body_y\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10606__X _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_330_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13622__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout208_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17269__A1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11002__A1 game.CPU.applesa.ab.absxs.body_x\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_326_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_303_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09746__A2 game.CPU.applesa.ab.check_walls.above.walls\[67\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11002__B2 game.CPU.applesa.ab.absxs.body_y\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09984_ game.CPU.apple_location2\[7\] _04208_ _04209_ net1489 vssd1 vssd1 vccd1 vccd1
+ _01380_ sky130_fd_sc_hd__a22o_1
XANTENNA__10761__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_243_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_271_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_243_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout744_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10501__B _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15580__A game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13463__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout532_X net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout911_A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18935__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09682__A1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1274_X net1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09682__B2 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_326_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09418_ net1146 game.CPU.applesa.ab.absxs.body_y\[97\] vssd1 vssd1 vccd1 vccd1 _03661_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10690_ _04592_ _04600_ _04672_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__o21a_1
XFILLER_0_325_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16952__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12428__B net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13766__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11332__B net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09434__A1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09349_ net926 game.CPU.applesa.ab.absxs.body_x\[11\] _03357_ net1159 _03591_ vssd1
+ vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__a221o_1
XFILLER_0_341_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09434__B2 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12360_ game.CPU.applesa.ab.absxs.body_x\[46\] net372 vssd1 vssd1 vccd1 vccd1 _06237_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_164_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16704__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15739__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11311_ game.CPU.applesa.ab.check_walls.above.walls\[65\] net772 vssd1 vssd1 vccd1
+ vccd1 _05200_ sky130_fd_sc_hd__xor2_1
X_12291_ game.CPU.applesa.ab.check_walls.above.walls\[14\] net419 vssd1 vssd1 vccd1
+ vccd1 _06177_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_321_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14030_ net959 _03468_ net787 net852 vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11242_ _03324_ net536 vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_238_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_276_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15755__A game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11173_ _03236_ net321 vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09753__A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ net1263 net1462 net1412 vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15981_ game.CPU.applesa.ab.check_walls.above.walls\[64\] net355 vssd1 vssd1 vccd1
+ vccd1 _01993_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_246_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_274_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_182_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17720_ _03085_ _03089_ _03090_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__nor3_1
XANTENNA__16289__C net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10055_ game.CPU.applesa.twoapples.count_luck\[4\] game.CPU.applesa.twoapples.count_luck\[3\]
+ _04261_ _04260_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__a31o_1
X_14932_ _08701_ _08708_ vssd1 vssd1 vccd1 vccd1 _08709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_215_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_261_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09903__D _04145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19710__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__B1 game.CPU.applesa.ab.check_walls.above.walls\[35\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17651_ _03037_ _03045_ _03046_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__and3_1
XANTENNA__11507__B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14863_ _08651_ net1787 vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[14\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_199_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16602_ net131 _02455_ net66 _02510_ game.writer.tracker.frame\[98\] vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.next_frame\[98\] sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_221_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13814_ _07684_ _07687_ net216 vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__mux2_1
X_17582_ game.CPU.kyle.L1.cnt_20ms\[5\] game.CPU.kyle.L1.cnt_20ms\[4\] _03002_ vssd1
+ vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__and3_1
XFILLER_0_202_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14794_ game.CPU.randy.counter1.count\[6\] _08608_ vssd1 vssd1 vccd1 vccd1 _08610_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19321_ clknet_leaf_70_clk _01345_ _00927_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.apple_location2_n\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_70_clk_X clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16533_ net113 _02468_ net716 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__o21a_1
XANTENNA__10807__A1 game.CPU.applesa.ab.absxs.body_y\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_329_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13745_ net246 _07590_ _07600_ _07618_ net180 vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__o311a_1
XFILLER_0_230_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10807__B2 game.CPU.applesa.ab.absxs.body_y\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17196__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10957_ _03287_ net412 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__nand2_1
XANTENNA__19860__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19252_ clknet_leaf_17_clk net1361 _00890_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_356_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16464_ net185 net117 _02418_ _02414_ net1873 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[56\]
+ sky130_fd_sc_hd__a32o_1
X_13676_ game.writer.tracker.frame\[494\] net841 net834 game.writer.tracker.frame\[493\]
+ vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__o22a_1
XANTENNA__16943__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10888_ net1172 net422 _04789_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__a21o_1
X_18203_ net580 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__inv_2
XANTENNA__12338__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13757__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15415_ _01428_ _01442_ game.writer.updater.commands.count\[15\] game.writer.updater.commands.count\[14\]
+ game.writer.updater.commands.count\[13\] vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_241_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11242__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12627_ game.CPU.applesa.ab.absxs.body_x\[59\] net530 net365 game.CPU.applesa.ab.absxs.body_y\[59\]
+ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19183_ clknet_leaf_5_clk _01302_ _00845_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_16395_ net245 _02367_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__or2_4
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_331_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18134_ net583 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_310_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15346_ game.writer.updater.commands.count\[2\] _08886_ game.writer.updater.commands.count\[4\]
+ game.writer.updater.commands.count\[3\] vssd1 vssd1 vccd1 vccd1 _08888_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12558_ game.CPU.applesa.ab.absxs.body_x\[85\] net375 net528 game.CPU.applesa.ab.absxs.body_x\[87\]
+ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_324_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12980__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18065_ net642 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11509_ _05397_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_232_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15277_ _01265_ _08827_ vssd1 vssd1 vccd1 vccd1 _08831_ sky130_fd_sc_hd__nor2_1
XANTENNA__12354__A game.CPU.applesa.ab.absxs.body_x\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold107 game.CPU.clock1.counter\[7\] vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ game.CPU.applesa.ab.absxs.body_x\[80\] net381 vssd1 vssd1 vccd1 vccd1 _06366_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_312_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold118 game.writer.tracker.frame\[372\] vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 game.writer.tracker.frame\[436\] vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_312_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17016_ _02509_ net86 net717 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__o21a_1
XFILLER_0_312_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14228_ game.CPU.applesa.ab.absxs.body_x\[41\] net1064 vssd1 vssd1 vccd1 vccd1 _08102_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_123_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_269_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19240__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_297_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14159_ net1104 net883 net944 net908 vssd1 vssd1 vccd1 vccd1 _08033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_284_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout609 net610 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_2
XFILLER_0_265_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09663__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18749__Q game.CPU.applesa.ab.absxs.body_x\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13288__A2 _07072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18967_ net1199 _00121_ _00638_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_23_clk_X clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_321_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ net604 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__inv_2
X_18898_ clknet_leaf_2_clk _00003_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA__19390__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1180 net1181 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_2
Xfanout1191 net1192 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__buf_2
X_17849_ _03173_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__inv_2
XANTENNA__17423__B2 net1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11417__B net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13445__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clk_X clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19519_ clknet_leaf_20_clk game.writer.tracker.next_frame\[114\] net1317 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[114\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_293_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout158_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16529__A3 _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13124__S net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_308_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_235_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11471__A1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_307_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12248__B net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09203_ game.CPU.applesa.ab.check_walls.above.walls\[138\] vssd1 vssd1 vccd1 vccd1
+ _03452_ sky130_fd_sc_hd__inv_2
XANTENNA__15654__A2_N net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_323_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12816__X _06690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout325_A net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10049__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_332_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1067_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ game.CPU.applesa.ab.check_walls.above.walls\[9\] vssd1 vssd1 vccd1 vccd1
+ _03383_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12420__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10991__B net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14463__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10577__A3 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09065_ game.CPU.applesa.ab.absxs.body_y\[31\] vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout113_X net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1234_A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 game.CPU.applesa.ab.count_luck\[5\] vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold641 game.writer.tracker.frame\[424\] vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout694_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold652 game.CPU.kyle.L1.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 game.writer.tracker.frame\[568\] vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1022_X net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_246_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10734__B1 _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19733__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09573__A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18659__Q game.CPU.applesa.ab.absxs.body_y\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout861_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ game.CPU.bodymain1.Direction\[0\] _04190_ vssd1 vssd1 vccd1 vccd1 _04196_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14476__A1 game.CPU.applesa.ab.absxs.body_x\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout959_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09292__B game.CPU.applesa.ab.check_walls.above.walls\[82\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09898_ _03819_ _03825_ _04139_ _04140_ _03577_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__o2111a_1
XANTENNA__09352__B1 game.CPU.applesa.ab.absxs.body_y\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13382__X _07256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19883__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16837__C net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ _05493_ _05745_ _05746_ _05747_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__and4_1
XFILLER_0_212_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10811_ net936 game.CPU.applesa.ab.absxs.body_y\[115\] net233 _04729_ vssd1 vssd1
+ vccd1 vccd1 _00986_ sky130_fd_sc_hd__a31o_1
X_11791_ _05673_ _05674_ _05677_ _05678_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_49_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09655__A1 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout914_X net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09655__B2 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_345_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_257_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13530_ _07402_ _07403_ net490 vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10742_ game.CPU.applesa.ab.absxs.body_y\[106\] _04658_ vssd1 vssd1 vccd1 vccd1 _04716_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_342_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_270_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16853__B _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11062__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13461_ net495 _07053_ net704 vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__a21o_1
X_10673_ net935 game.CPU.applesa.ab.absxs.body_x\[115\] net233 _04703_ vssd1 vssd1
+ vccd1 vccd1 _01098_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_341_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_313_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15200_ _03524_ game.CPU.applesa.normal1.number\[0\] game.CPU.applesa.normal1.number\[1\]
+ vssd1 vssd1 vccd1 vccd1 _08769_ sky130_fd_sc_hd__o21ai_1
XANTENNA__16572__C net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_298_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12412_ game.CPU.applesa.ab.absxs.body_x\[55\] net532 net365 game.CPU.applesa.ab.absxs.body_y\[55\]
+ _06288_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__a221o_1
XANTENNA__12411__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16180_ _01758_ _01763_ _02160_ _02191_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__or4_1
X_13392_ net697 _06891_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__or2_1
XANTENNA__19263__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15131_ net1208 net1233 net788 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__and3_1
XANTENNA__17965__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12343_ _03244_ net374 vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16153__B2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_346_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12274_ game.CPU.applesa.ab.check_walls.above.walls\[158\] net418 vssd1 vssd1 vccd1
+ vccd1 _06160_ sky130_fd_sc_hd__xnor2_1
X_15062_ net1218 net1247 game.CPU.applesa.ab.check_walls.above.walls\[90\] vssd1 vssd1
+ vccd1 vccd1 _00285_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11517__A2 _05210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_268_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11225_ game.CPU.applesa.ab.absxs.body_y\[12\] net535 vssd1 vssd1 vccd1 vccd1 _05115_
+ sky130_fd_sc_hd__or2_1
XANTENNA__13911__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14013_ net938 net781 vssd1 vssd1 vccd1 vccd1 _07887_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_130_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19870_ clknet_leaf_27_clk game.writer.tracker.next_frame\[465\] net1311 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[465\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09591__B1 game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18821_ clknet_leaf_2_clk _01212_ vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dfxtp_1
X_11156_ _03271_ net544 vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__nand2_1
XANTENNA__18569__Q game.CPU.applesa.ab.absxs.body_y\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_262_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_235_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15664__B1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_297_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10107_ _04313_ net1489 _04311_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__mux2_1
X_18752_ clknet_leaf_59_clk _01169_ _00489_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[38\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11518__A _03380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11087_ _03305_ net539 vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__nand2_1
X_15964_ _01966_ _01967_ _01974_ _01975_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__or4_2
XANTENNA__12478__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17703_ _03076_ _03077_ _03080_ vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__and3_1
XFILLER_0_222_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10038_ _04210_ _04212_ _04224_ _04232_ game.CPU.applesa.twoapples.collisions vssd1
+ vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__a41o_1
X_14915_ _08424_ _08426_ _08428_ _08430_ vssd1 vssd1 vccd1 vccd1 _08692_ sky130_fd_sc_hd__and4_1
XANTENNA__15932__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18683_ clknet_leaf_8_clk _01100_ _00420_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_15895_ game.CPU.applesa.ab.absxs.body_y\[43\] net436 vssd1 vssd1 vccd1 vccd1 _01907_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_349_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13690__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16759__A3 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_357_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ _08811_ _03009_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__nor2_1
X_14846_ net1691 _08641_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[7\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_187_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17565_ _02783_ _02839_ net426 vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__a21oi_1
X_14777_ _08586_ _08590_ _08597_ vssd1 vssd1 vccd1 vccd1 _08598_ sky130_fd_sc_hd__nor3_1
XANTENNA__09646__A1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_141_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_336_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09646__B2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ game.CPU.applesa.ab.check_walls.above.walls\[182\] net290 net296 game.CPU.applesa.ab.check_walls.above.walls\[183\]
+ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a2bb2o_1
X_19304_ clknet_leaf_56_clk game.CPU.applesa.ab.check_walls.collision_rightn _00919_
+ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.collision_right sky130_fd_sc_hd__dfrtp_1
X_16516_ _02267_ net152 vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__and2_2
X_13728_ game.writer.tracker.frame\[249\] game.writer.tracker.frame\[251\] game.writer.tracker.frame\[252\]
+ game.writer.tracker.frame\[250\] net981 net1031 vssd1 vssd1 vccd1 vccd1 _07602_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17496_ net1258 _02843_ _02924_ net1274 _02829_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__a32o_1
XFILLER_0_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11453__B2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_50_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17184__A3 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19235_ clknet_leaf_7_clk _00066_ _00873_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_16447_ net238 net236 _02296_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__or3_4
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19606__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13659_ game.writer.tracker.frame\[41\] game.writer.tracker.frame\[43\] game.writer.tracker.frame\[44\]
+ game.writer.tracker.frame\[42\] net970 net992 vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__mux4_1
XFILLER_0_305_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14564__A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19166_ clknet_leaf_57_clk _01286_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count_luck\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16378_ net172 _02289_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__nand2_2
XFILLER_0_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12953__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18117_ net582 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11700__B net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15329_ _00029_ _08869_ _08870_ _08871_ _08872_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__o32a_1
XFILLER_0_124_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09377__B net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19097_ net1178 _00135_ _00768_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[142\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_65_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16144__A1 game.CPU.applesa.ab.absxs.body_x\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12084__A game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15098__C net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16144__B2 game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_41_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18630__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19756__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18048_ net660 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_312_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13908__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__B1 _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout406 net407 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_4
XFILLER_0_39_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20010_ net1379 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout417 net418 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09821_ _04058_ _04059_ _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__or3_2
Xfanout428 _02818_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_2
Xfanout439 _08429_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_4
X_19999_ clknet_leaf_44_clk _01423_ net1299 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_226_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16003__B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18780__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11428__A game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09752_ net1160 net826 vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__nand2_1
XANTENNA__12469__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13666__C1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Left_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_280_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15842__B net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09683_ net899 game.CPU.applesa.ab.absxs.body_y\[101\] _03921_ _03924_ _03925_ vssd1
+ vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout275_A _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_241_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_275_Right_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19136__CLK net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11692__A1 game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13418__C1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14458__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10986__B net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_355_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout442_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19103__Q game.CPU.applesa.ab.check_walls.above.walls\[148\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12259__A game.CPU.applesa.ab.check_walls.above.walls\[165\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1184_A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_18_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16907__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_308_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16673__B net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13789__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout57 _02692_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_2
XANTENNA__19286__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout230_X net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout68 _02373_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1351_A net1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_312_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout79 net82 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_2
XFILLER_0_134_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13816__S0 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_114_Left_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13197__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_312_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14193__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12944__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ game.writer.updater.commands.cmd_num\[2\] vssd1 vssd1 vccd1 vccd1 _03366_
+ sky130_fd_sc_hd__inv_2
XANTENNA__09287__B game.CPU.applesa.ab.check_walls.above.walls\[83\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10507__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1237_X net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_304_Left_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_288_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12604__A2_N net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09048_ game.CPU.applesa.ab.absxs.body_y\[93\] vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__inv_2
XANTENNA__14146__B1 _08017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19773__Q game.writer.tracker.frame\[368\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold460 game.writer.tracker.frame\[211\] vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12722__A _06571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout90_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold471 game.CPU.walls.rand_wall.count_luck\[7\] vssd1 vssd1 vccd1 vccd1 net1856
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 game.writer.tracker.frame\[377\] vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ game.CPU.applesa.ab.absxs.body_y\[55\] net398 vssd1 vssd1 vccd1 vccd1 _04900_
+ sky130_fd_sc_hd__xnor2_1
Xhold493 game.writer.tracker.frame\[260\] vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout940 game.CPU.applesa.y\[3\] vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_123_Left_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11338__A game.CPU.applesa.ab.check_walls.above.walls\[81\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout951 net957 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_8
Xfanout962 net963 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__buf_4
Xfanout973 net982 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_2
Xfanout984 net1042 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_8
Xfanout995 net997 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_273_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12961_ net513 _06834_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__or2_1
XANTENNA__15752__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14700_ game.CPU.randy.counter1.count1\[11\] _08491_ _08514_ _08538_ vssd1 vssd1
+ vccd1 vccd1 _08539_ sky130_fd_sc_hd__a211o_1
XANTENNA__16567__C _02415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_313_Left_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09750__B game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11912_ game.CPU.applesa.ab.check_walls.above.walls\[12\] net393 net302 game.CPU.applesa.ab.check_walls.above.walls\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__o22ai_1
XPHY_EDGE_ROW_242_Right_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15680_ game.CPU.applesa.ab.check_walls.above.walls\[14\] net442 vssd1 vssd1 vccd1
+ vccd1 _01692_ sky130_fd_sc_hd__nor2_1
XANTENNA__10486__A2 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12892_ _06762_ _06763_ _06764_ _06765_ net497 net690 vssd1 vssd1 vccd1 vccd1 _06766_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_358_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14368__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14631_ game.CPU.clock1.counter\[16\] _08475_ net267 vssd1 vssd1 vccd1 vccd1 _08477_
+ sky130_fd_sc_hd__o21ai_1
X_11843_ _05721_ _05722_ _05730_ net192 vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__a31o_1
XFILLER_0_353_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19629__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12176__A1_N net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17350_ _02773_ _02779_ _02777_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__o21ai_1
X_14562_ game.CPU.walls.abc.enable game.CPU.walls.abc.number_out\[6\] vssd1 vssd1
+ vccd1 vccd1 _08428_ sky130_fd_sc_hd__nand2_2
XANTENNA__12632__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11774_ net793 net390 _05657_ _05658_ _05661_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_132_Left_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17166__A3 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16301_ _02273_ _02300_ _02293_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[11\]
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_103_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ net683 _07126_ _07365_ net209 vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__o211a_1
X_17281_ net117 _02576_ _02751_ net1936 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[540\]
+ sky130_fd_sc_hd__a22o_1
X_10725_ game.CPU.applesa.ab.absxs.body_y\[37\] _04642_ _04643_ game.CPU.applesa.ab.absxs.body_y\[33\]
+ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_222_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14493_ _08275_ _08279_ _08164_ _08173_ _08196_ vssd1 vssd1 vccd1 vccd1 _08367_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19020_ net1202 _00249_ _00691_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[65\]
+ sky130_fd_sc_hd__dfrtp_4
X_16232_ net141 _02239_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__or2_4
XANTENNA__18653__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_190_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09478__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13444_ _06932_ _06938_ net682 vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__mux2_1
XANTENNA__19779__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10656_ game.CPU.applesa.ab.absxs.body_x\[34\] _04696_ _04697_ game.CPU.applesa.ab.absxs.body_x\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11199__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12616__B _06492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_322_Left_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17695__A game.CPU.walls.rand_wall.input2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16163_ _02071_ _02078_ _02174_ _02150_ _01963_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__o311a_1
XANTENNA__11520__B net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload16 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload16/X sky130_fd_sc_hd__clkbuf_4
X_13375_ _06658_ _06696_ _06698_ _06699_ net502 net694 vssd1 vssd1 vccd1 vccd1 _07249_
+ sky130_fd_sc_hd__mux4_1
X_10587_ net1080 _04665_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__nor2_2
Xclkload27 clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__inv_12
Xclkload38 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__09800__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload49 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload49/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09800__B2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_279_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15114_ net1204 net1231 net791 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__and3_1
X_12326_ net375 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.absxs.next_head\[1\]
+ sky130_fd_sc_hd__inv_4
X_16094_ game.CPU.applesa.ab.absxs.body_y\[109\] net337 vssd1 vssd1 vccd1 vccd1 _02106_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19009__CLK net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13287__X _07161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19922_ clknet_leaf_33_clk game.writer.tracker.next_frame\[517\] net1302 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[517\] sky130_fd_sc_hd__dfrtp_1
X_15045_ net1217 net1244 game.CPU.applesa.ab.check_walls.above.walls\[73\] vssd1 vssd1
+ vccd1 vccd1 _00267_ sky130_fd_sc_hd__and3_1
X_12257_ net822 net419 vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_71_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11208_ _03297_ net405 vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__xnor2_1
X_19853_ clknet_leaf_36_clk game.writer.tracker.next_frame\[448\] net1356 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[448\] sky130_fd_sc_hd__dfrtp_1
X_12188_ _05955_ _05956_ _06072_ _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__or4_1
XANTENNA__16598__X _02512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12351__B net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11910__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18804_ clknet_leaf_1_clk game.CPU.clock1.next_counter\[7\] _00541_ vssd1 vssd1 vccd1
+ vccd1 game.CPU.clock1.counter\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_305_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11139_ _05019_ _05021_ _05024_ _05027_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__or4_1
XANTENNA__19159__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19784_ clknet_leaf_23_clk game.writer.tracker.next_frame\[379\] net1347 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[379\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13648__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16996_ _02566_ net85 net558 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_262_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_331_Left_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18735_ clknet_leaf_16_clk _01152_ _00472_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[105\]
+ sky130_fd_sc_hd__dfrtp_4
X_15947_ game.CPU.applesa.ab.check_walls.above.walls\[42\] net469 vssd1 vssd1 vccd1
+ vccd1 _01959_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18666_ clknet_leaf_70_clk _01083_ _00403_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[92\]
+ sky130_fd_sc_hd__dfrtp_4
X_15878_ _01881_ _01885_ _01888_ _01889_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__or4_1
X_17617_ game.CPU.kyle.L1.cnt_20ms\[11\] game.CPU.kyle.L1.cnt_20ms\[10\] _03023_ vssd1
+ vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_69_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14829_ game.CPU.randy.f1.c1.count\[0\] game.CPU.randy.f1.c1.count\[1\] _08631_ vssd1
+ vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[1\] sky130_fd_sc_hd__o21a_1
X_18597_ clknet_leaf_60_clk _01017_ _00334_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[74\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_263_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17548_ _04484_ _02837_ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_290_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16493__B net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17479_ _02905_ _02907_ _02904_ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13402__S net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19218_ clknet_leaf_68_clk _01312_ _00857_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_location\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_154_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17101__C net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12526__B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12926__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19149_ net1187 _00192_ _00820_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[194\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11430__B net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17314__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10937__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14128__B1 game.CPU.applesa.ab.check_walls.above.walls\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15837__B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15876__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_344_Right_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13964__A2_N game.CPU.applesa.ab.check_walls.above.walls\[177\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16014__A game.CPU.applesa.ab.check_walls.above.walls\[176\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13351__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout203 net208 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_4
Xfanout214 net217 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_243_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout225 net232 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout392_A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12261__B net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11362__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 net237 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout247 net248 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_4
XANTENNA__13925__X _07799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09804_ _04043_ _04044_ _04045_ _04046_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__or4_1
XANTENNA__15853__A game.CPU.applesa.ab.absxs.body_y\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11158__A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout258 _05195_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_4
Xfanout269 game.CPU.walls.rand_wall.abduyd.next_wall\[0\] vssd1 vssd1 vccd1 vccd1
+ net269 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16668__B net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09851__A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16840__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09735_ net915 game.CPU.applesa.ab.absxs.body_x\[33\] game.CPU.applesa.ab.absxs.body_y\[35\]
+ net907 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout657_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10468__A2 game.CPU.applesa.ab.absxs.body_x\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09666_ _03906_ _03907_ _03908_ _03905_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__a211o_1
XANTENNA__16053__B1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09597_ net1109 game.CPU.applesa.ab.absxs.body_x\[72\] vssd1 vssd1 vccd1 vccd1 _03840_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__09997__S _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15800__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18676__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_254_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19921__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18672__Q game.CPU.applesa.ab.absxs.body_y\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_176_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10510_ game.CPU.applesa.ab.absxs.body_x\[69\] _04625_ _04626_ game.CPU.applesa.ab.absxs.body_x\[65\]
+ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__a22o_1
XANTENNA__09298__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11490_ _05378_ _05249_ _05234_ _05217_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_118_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_351_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12436__B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16825__A_N _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10441_ net1438 net849 _04171_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__a21o_1
XFILLER_0_162_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16108__B2 game.CPU.applesa.ab.absxs.body_y\[38\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_162_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10928__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16659__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16850__C net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12393__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13160_ game.writer.tracker.frame\[158\] game.writer.tracker.frame\[159\] net1023
+ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__mux2_1
X_10372_ net1445 net848 _04203_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout981_X net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15747__B net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_343_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12111_ game.CPU.applesa.ab.check_walls.above.walls\[52\] net553 vssd1 vssd1 vccd1
+ vccd1 _05998_ sky130_fd_sc_hd__nand2_1
X_13091_ game.writer.tracker.frame\[238\] game.writer.tracker.frame\[239\] net998
+ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__mux2_1
XANTENNA__12452__A game.CPU.applesa.ab.absxs.body_y\[50\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_311_Right_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_265_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12042_ _05476_ _05480_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_236_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold290 game.writer.tracker.frame\[363\] vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_207_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_291_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19008__Q game.CPU.applesa.ab.check_walls.above.walls\[53\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17084__A2 _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16850_ net131 net67 net143 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__and3_1
XFILLER_0_217_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout770 net772 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__clkbuf_8
X_15801_ _01806_ _01811_ _01812_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__and3_1
Xfanout781 game.CPU.applesa.ab.check_walls.above.walls\[191\] vssd1 vssd1 vccd1 vccd1
+ net781 sky130_fd_sc_hd__clkbuf_4
X_16781_ net152 _02454_ net107 _02595_ net1641 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[196\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_189_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout792 game.CPU.applesa.ab.check_walls.above.walls\[133\] vssd1 vssd1 vccd1 vccd1
+ net792 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09849__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13993_ net1061 game.CPU.applesa.ab.check_walls.above.walls\[73\] vssd1 vssd1 vccd1
+ vccd1 _07867_ sky130_fd_sc_hd__xor2_1
XANTENNA__13645__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09849__B2 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18520_ net581 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15732_ game.CPU.applesa.ab.absxs.body_y\[12\] net452 vssd1 vssd1 vccd1 vccd1 _01744_
+ sky130_fd_sc_hd__xnor2_1
X_12944_ net200 _06739_ _06817_ net282 vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__a211o_1
XANTENNA__16044__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_354_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ net652 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
XFILLER_0_358_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15663_ net436 game.CPU.applesa.ab.check_walls.above.walls\[55\] _03406_ net352 vssd1
+ vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__16595__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ game.writer.tracker.frame\[2\] game.writer.tracker.frame\[4\] game.writer.tracker.frame\[5\]
+ game.writer.tracker.frame\[3\] net969 net1002 vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__mux4_1
XANTENNA__16594__A _02351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17402_ net1264 game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__nand2_1
X_14614_ _08465_ _08466_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[9\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_276_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12605__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18382_ net600 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__inv_2
X_11826_ game.CPU.applesa.ab.check_walls.above.walls\[125\] net305 vssd1 vssd1 vccd1
+ vccd1 _05714_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15594_ game.CPU.applesa.ab.check_walls.above.walls\[37\] net338 vssd1 vssd1 vccd1
+ vccd1 _01606_ sky130_fd_sc_hd__nand2_1
XANTENNA__19678__Q game.writer.tracker.frame\[273\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17139__A3 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_218_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17333_ _01440_ _01579_ _02765_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a21o_1
XFILLER_0_157_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16347__A1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14545_ net356 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.abduyd.next_wall\[0\]
+ sky130_fd_sc_hd__clkinv_4
XFILLER_0_327_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11757_ net783 net311 vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17264_ net162 net70 _02479_ net724 vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__o31a_1
XANTENNA__16898__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10708_ net1270 net425 _04710_ net933 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__a22o_1
XFILLER_0_342_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14476_ game.CPU.applesa.ab.absxs.body_x\[9\] net883 net1050 _03289_ vssd1 vssd1
+ vccd1 vccd1 _08350_ sky130_fd_sc_hd__o22a_1
XANTENNA__10418__Y _04563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11688_ game.CPU.applesa.ab.check_walls.above.walls\[61\] net317 vssd1 vssd1 vccd1
+ vccd1 _05577_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12346__B net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19003_ net1195 _00230_ _00674_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[48\]
+ sky130_fd_sc_hd__dfrtp_4
X_16215_ _06571_ net835 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__nor2_2
X_13427_ _06944_ _06946_ net702 vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17195_ _02503_ net74 _02729_ net1546 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[476\]
+ sky130_fd_sc_hd__a22o_1
X_10639_ net932 game.CPU.applesa.ab.absxs.body_x\[45\] net561 _04687_ vssd1 vssd1
+ vccd1 vccd1 _01116_ sky130_fd_sc_hd__a31o_1
XANTENNA_max_cap455_A net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18314__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16146_ _03436_ net270 vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09936__A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13358_ _06662_ _06664_ net703 vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15657__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_307_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12309_ game.CPU.applesa.ab.check_walls.above.walls\[190\] net418 vssd1 vssd1 vccd1
+ vccd1 _06195_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_287_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16077_ _03231_ net343 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__xnor2_1
X_13289_ _07047_ _07162_ net174 vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_219_Left_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12362__A game.CPU.applesa.ab.absxs.body_x\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13333__A1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19905_ clknet_leaf_20_clk game.writer.tracker.next_frame\[500\] net1316 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[500\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_229_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15028_ net1222 net1256 game.CPU.applesa.ab.check_walls.above.walls\[56\] vssd1 vssd1
+ vccd1 vccd1 _00248_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17075__A2 net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15673__A game.CPU.applesa.ab.check_walls.above.walls\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_19836_ clknet_leaf_33_clk game.writer.tracker.next_frame\[431\] net1325 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[431\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10698__A2 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16121__X _02133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16822__A2 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_223_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18757__Q game.CPU.applesa.ab.absxs.body_x\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13097__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19767_ clknet_leaf_28_clk game.writer.tracker.next_frame\[362\] net1288 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[362\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13905__B game.CPU.applesa.ab.check_walls.above.walls\[120\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16979_ net152 _02454_ net90 _02665_ net1556 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[324\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__13636__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 gpio_in[1] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09520_ _03759_ _03760_ _03761_ _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__a22o_1
XANTENNA__09390__B net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18718_ clknet_leaf_70_clk _01135_ _00455_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[88\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__18699__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19698_ clknet_leaf_29_clk game.writer.tracker.next_frame\[293\] net1284 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[293\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19944__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09451_ _03685_ _03689_ _03693_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_318_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18649_ clknet_leaf_12_clk _01066_ _00386_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[55\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_228_Left_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_160_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14597__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09382_ net1103 _03383_ game.CPU.applesa.ab.check_walls.above.walls\[14\] net904
+ _03624_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__a221o_1
XFILLER_0_337_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13495__S1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13132__S net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16889__A2 _02456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10622__A2 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11160__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout405_A game.CPU.applesa.ab.absxs.next_head\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18224__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1147_A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16670__C net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09776__B1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09846__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_329_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_237_Left_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09565__B game.CPU.applesa.ab.absxs.body_x\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12272__A game.CPU.applesa.ab.check_walls.above.walls\[157\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1314_A net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1009 net1042 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout774_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19474__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16679__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_273_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1102_X net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16398__B _02280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16813__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout941_A game.CPU.applesa.y\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13183__S0 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_260_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09718_ net1126 game.CPU.applesa.ab.absxs.body_y\[87\] vssd1 vssd1 vccd1 vccd1 _03961_
+ sky130_fd_sc_hd__or2_1
X_10990_ game.CPU.applesa.ab.absxs.body_y\[115\] net398 vssd1 vssd1 vccd1 vccd1 _04880_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout53_A _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_241_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09700__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09649_ _03886_ _03891_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__or2_4
XFILLER_0_328_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_355_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11845__A1_N game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12660_ game.CPU.applesa.ab.absxs.body_x\[67\] net532 net521 game.CPU.applesa.ab.absxs.body_y\[66\]
+ _06375_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__a221o_1
XFILLER_0_328_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11611_ net803 net257 vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__or2_1
XFILLER_0_167_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12591_ game.CPU.applesa.ab.absxs.body_x\[58\] net373 vssd1 vssd1 vccd1 vccd1 _06468_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_100_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13042__S net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14330_ _03267_ net1063 net962 _03332_ vssd1 vssd1 vccd1 vccd1 _08204_ sky130_fd_sc_hd__o22a_1
X_11542_ net773 _05430_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11810__A1 game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12166__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_279_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14261_ _08132_ _08133_ _08134_ _08131_ vssd1 vssd1 vccd1 vccd1 _08135_ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12881__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15552__A2 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire456 _08425_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_2
X_11473_ net818 net261 vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__or2_1
X_16000_ _03431_ net270 net439 net803 _02011_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__o221a_1
X_13212_ net214 _07077_ _07085_ net279 vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__a211o_1
XANTENNA__13563__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_213_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10424_ _04567_ _04568_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__nand2_1
X_14192_ _03261_ net1061 net1045 _03260_ vssd1 vssd1 vccd1 vccd1 _08066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19817__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13143_ game.writer.tracker.frame\[146\] game.writer.tracker.frame\[147\] net1023
+ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16501__A1 _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10355_ net2032 _04516_ _04520_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12182__A game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13315__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14512__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13074_ game.writer.tracker.frame\[232\] game.writer.tracker.frame\[233\] net998
+ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__mux2_1
X_10286_ net851 game.CPU.applesa.ab.y_final\[1\] game.CPU.applesa.ab.good_spot_next
+ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__and3_1
X_17951_ net607 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_295_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17057__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16902_ _02309_ net92 _02642_ net1630 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[270\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_228_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12025_ net829 net297 vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__xnor2_1
X_17882_ net637 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__inv_2
X_19621_ clknet_leaf_21_clk game.writer.tracker.next_frame\[216\] net1336 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[216\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19967__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18577__Q game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_302_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16833_ _02525_ net98 net715 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__o21a_1
XANTENNA__16101__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11526__A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16764_ net185 _02418_ net109 _02590_ net1632 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[184\]
+ sky130_fd_sc_hd__a32o_1
X_19552_ clknet_leaf_34_clk game.writer.tracker.next_frame\[147\] net1319 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[147\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_205_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13976_ net868 net810 game.CPU.applesa.ab.check_walls.above.walls\[85\] net862 vssd1
+ vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__a22o_1
XFILLER_0_232_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18503_ net587 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__inv_2
XANTENNA_output34_A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15715_ _03291_ net351 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__xnor2_1
X_12927_ _06682_ _06689_ net220 vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__mux2_1
XANTENNA__15940__B net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19483_ clknet_leaf_18_clk game.writer.tracker.next_frame\[78\] net1308 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[78\] sky130_fd_sc_hd__dfrtp_1
X_16695_ _02311_ net61 net556 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12909__X _06783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16568__B2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_200_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18434_ net581 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15646_ _03422_ net456 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__xnor2_1
X_12858_ game.writer.tracker.frame\[298\] game.writer.tracker.frame\[299\] net988
+ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_346_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18365_ net596 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__inv_2
XANTENNA__12054__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11809_ net817 net393 _05693_ _05571_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_196_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12054__B2 game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15577_ game.CPU.applesa.ab.check_walls.above.walls\[90\] net469 vssd1 vssd1 vccd1
+ vccd1 _01589_ sky130_fd_sc_hd__xnor2_1
X_12789_ game.writer.tracker.frame\[384\] game.writer.tracker.frame\[385\] net1032
+ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_346_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12357__A game.CPU.applesa.ab.absxs.body_x\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_346_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17316_ net1743 _02761_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[565\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_56_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14528_ _07400_ _08370_ vssd1 vssd1 vccd1 vccd1 _08402_ sky130_fd_sc_hd__or2_1
XANTENNA__19347__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10604__A2 _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18296_ net620 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_313_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17247_ net111 _02452_ _02742_ net1569 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[515\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14459_ _03251_ net1067 net964 _03319_ _08324_ vssd1 vssd1 vccd1 vccd1 _08333_ sky130_fd_sc_hd__a221o_1
XANTENNA__16740__A1 _02375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12644__X _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17178_ _02476_ net73 _02725_ net1874 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[463\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10368__A1 game.CPU.applesa.ab.absxs.body_y\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14291__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19497__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16129_ _01663_ _01665_ _02137_ _02138_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__or4_1
XFILLER_0_141_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_330_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19962__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17296__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14503__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08951_ net1144 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11317__B1 game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17048__A2 _02412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13916__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_324_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11014__A2_N net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19819_ clknet_leaf_38_clk game.writer.tracker.next_frame\[414\] net1333 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[414\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_208_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_162_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10540__A1 _03197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16011__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13165__S0 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13127__S net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout188_A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09503_ net1101 _03406_ game.CPU.applesa.ab.check_walls.above.walls\[50\] net922
+ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11155__B net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_338_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15850__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13490__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout355_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_296_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1097_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17220__A2 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ net1131 _03337_ _03338_ net1141 _03676_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10994__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_304_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09365_ _03600_ _03606_ _03607_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout143_X net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19111__Q game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout522_A _06214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_325_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_30 _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ _03537_ _03538_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_41 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_52 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_340_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18714__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15578__A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_245_Left_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16731__A1 _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1052_X net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout891_A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout989_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17287__A2 _02512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_249_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16495__B1 _02357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10140_ game.CPU.randy.f1.a1.count\[11\] game.CPU.randy.f1.a1.count\[10\] game.CPU.randy.f1.a1.count\[9\]
+ game.CPU.randy.f1.a1.count\[8\] vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_329_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_274_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19781__Q game.writer.tracker.frame\[376\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_262_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13848__A2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17039__A2 _02391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ _04272_ _04278_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__and2b_1
XANTENNA__11859__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17444__C1 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_254_Left_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13830_ game.writer.tracker.frame\[543\] net708 net835 game.writer.tracker.frame\[541\]
+ net507 vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__o221a_1
XANTENNA__12808__A0 _06678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout56_X net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11065__B net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13761_ net482 _07633_ _07634_ vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__and3_1
XANTENNA__15760__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13481__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973_ game.CPU.applesa.ab.absxs.body_y\[75\] net397 vssd1 vssd1 vccd1 vccd1 _04863_
+ sky130_fd_sc_hd__nor2_1
X_15500_ net870 net853 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17211__A2 _02375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13561__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12712_ _06585_ _06584_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__and2b_1
X_16480_ net1837 _02426_ _02429_ net112 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[61\]
+ sky130_fd_sc_hd__a22o_1
X_13692_ game.writer.tracker.frame\[507\] net710 net673 game.writer.tracker.frame\[508\]
+ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14376__B net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_273_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15431_ _01440_ _01458_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__or2_1
XFILLER_0_214_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17968__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12643_ _06259_ _06449_ _06450_ _06519_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__or4_1
XANTENNA__16970__A1 _02435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19021__Q game.CPU.applesa.ab.check_walls.above.walls\[66\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_343_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18150_ net630 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15362_ _08903_ vssd1 vssd1 vccd1 vccd1 _08904_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_263_Left_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12574_ game.CPU.applesa.ab.absxs.body_y\[5\] net526 net367 game.CPU.applesa.ab.absxs.body_y\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__o22a_1
X_17101_ net185 _02498_ net80 vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__and3_1
XANTENNA__10598__B2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14313_ game.CPU.applesa.ab.absxs.body_x\[58\] net1059 vssd1 vssd1 vccd1 vccd1 _08187_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_182_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18081_ net663 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ game.CPU.applesa.ab.check_walls.above.walls\[41\] net771 vssd1 vssd1 vccd1
+ vccd1 _05414_ sky130_fd_sc_hd__xor2_1
XFILLER_0_312_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15293_ _00029_ _08842_ vssd1 vssd1 vccd1 vccd1 _08843_ sky130_fd_sc_hd__nand2_1
XANTENNA__16722__B2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17032_ _02377_ _02678_ _02681_ net1861 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[361\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_349_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14244_ game.CPU.applesa.ab.absxs.body_x\[23\] net1046 vssd1 vssd1 vccd1 vccd1 _08118_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_230_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11456_ game.CPU.applesa.ab.check_walls.above.walls\[76\] net253 _05340_ _05341_
+ _05344_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_312_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17278__A2 _02258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10407_ game.CPU.randy.f1.state\[1\] _04341_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__or2_1
XANTENNA__15000__B net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14175_ _03254_ net1067 net874 game.CPU.applesa.ab.absxs.body_x\[107\] _08048_ vssd1
+ vssd1 vccd1 vccd1 _08049_ sky130_fd_sc_hd__a221o_1
X_11387_ _03479_ net257 vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13126_ net224 _06999_ _06992_ net274 vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_284_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10338_ _04490_ _04511_ game.CPU.randy.f1.a1.count\[6\] net739 vssd1 vssd1 vccd1
+ vccd1 _01296_ sky130_fd_sc_hd__a2bb2o_1
X_18983_ net1197 _00208_ _00654_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10770__A1 game.CPU.applesa.ab.absxs.body_y\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_226_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ game.writer.tracker.frame\[220\] game.writer.tracker.frame\[221\] net1016
+ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__mux2_1
X_17934_ net659 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_272_Left_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10269_ net759 net563 vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__or2_1
Xfanout1340 net1341 vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__buf_2
XFILLER_0_280_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12008_ net813 _05192_ _05863_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__and3_1
XANTENNA__12511__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1351 net1353 vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_252_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16789__A1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17865_ game.writer.updater.commands.count\[14\] game.writer.updater.commands.count\[13\]
+ _03180_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__and3_1
X_19604_ clknet_leaf_19_clk game.writer.tracker.next_frame\[199\] net1342 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[199\] sky130_fd_sc_hd__dfrtp_1
X_16816_ _02509_ net98 net727 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__o21a_1
X_17796_ net879 _03134_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14264__A2 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19535_ clknet_leaf_32_clk game.writer.tracker.next_frame\[130\] net1301 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[130\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_198_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15670__B net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16747_ _02390_ net101 _02583_ net1726 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[173\]
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_187_Right_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13959_ net939 net783 vssd1 vssd1 vccd1 vccd1 _07833_ sky130_fd_sc_hd__nand2_1
XANTENNA__14567__A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_242_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_315_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19466_ clknet_leaf_40_clk game.writer.tracker.next_frame\[61\] net1358 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[61\] sky130_fd_sc_hd__dfrtp_1
X_16678_ net174 _02237_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__nor2_1
XFILLER_0_319_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_335_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18417_ net627 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__inv_2
XANTENNA__18737__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15629_ game.CPU.applesa.ab.check_walls.above.walls\[184\] net354 net430 net781 vssd1
+ vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__16961__A1 _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_281_Left_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_271_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19397_ clknet_leaf_47_clk game.writer.control.next\[0\] net1298 vssd1 vssd1 vccd1
+ vccd1 game.writer.control.current\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12087__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13775__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09979__B1 _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ net824 vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__inv_2
X_18348_ net594 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10319__B net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12983__C1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09081_ game.CPU.applesa.ab.absxs.body_y\[81\] vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__inv_2
X_18279_ net644 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16713__A1 _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09396__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18887__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload42_A clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13622__S1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16006__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17269__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11002__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_326_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout103_A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09983_ _03518_ _04208_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__nor2_2
XANTENNA__15845__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11718__X _05606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__A game.CPU.applesa.ab.absxs.body_y\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1012_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10989__B net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout472_A net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19106__Q game.CPU.applesa.ab.check_walls.above.walls\[151\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13138__S0 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17441__A2 _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19512__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15580__B net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout260_X net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_337_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout737_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09417_ net1083 game.CPU.applesa.ab.absxs.body_x\[99\] vssd1 vssd1 vccd1 vccd1 _03660_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_338_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19662__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16952__A1 _02405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout904_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1267_X net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12569__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09348_ net1132 game.CPU.applesa.ab.absxs.body_y\[11\] vssd1 vssd1 vccd1 vccd1 _03591_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_325_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14483__Y _08357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_325_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16704__A1 _02322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ net757 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__inv_2
XANTENNA__12725__A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_340_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11310_ _05198_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12290_ _06175_ _05916_ _05914_ _06174_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_210_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11241_ game.CPU.applesa.ab.absxs.body_y\[109\] net542 vssd1 vssd1 vccd1 vccd1 _05131_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_132_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15755__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ _05058_ _05059_ _05060_ _05061_ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__a22o_1
XANTENNA__19042__CLK net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_289_Right_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_246_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10752__B2 game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10123_ game.CPU.applesa.ab.start_enable game.CPU.applesa.ab.good_collision vssd1
+ vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__or2_1
XFILLER_0_274_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09753__B net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15980_ game.CPU.applesa.ab.check_walls.above.walls\[71\] net434 vssd1 vssd1 vccd1
+ vccd1 _01992_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_234_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_262_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_261_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10054_ game.CPU.applesa.twoapples.count_luck\[4\] game.CPU.applesa.twoapples.count_luck\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__nand2_1
X_14931_ _08704_ _08707_ vssd1 vssd1 vccd1 vccd1 _08708_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10504__A1 game.CPU.applesa.ab.absxs.body_x\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_292_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19016__Q game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10504__B2 game.CPU.applesa.ab.absxs.body_x\[73\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09370__A1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17650_ game.CPU.kyle.L1.cnt_500hz\[7\] _03044_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__nand2_1
X_14862_ game.CPU.randy.f1.c1.count\[13\] _08649_ net1786 vssd1 vssd1 vccd1 vccd1
+ _08652_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09370__B2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19192__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16586__B _02387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13813_ _07685_ _07686_ net497 vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__mux2_1
X_16601_ _02447_ _02451_ net206 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_242_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_221_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ game.CPU.kyle.L1.cnt_20ms\[3\] _03001_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14793_ _08608_ _08609_ net138 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__and3b_1
XANTENNA__12459__X _06336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14387__A game.CPU.applesa.ab.absxs.body_y\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16532_ net159 _02303_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__or2_2
X_19320_ clknet_leaf_71_clk _01344_ _00926_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.apple_location2_n\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11804__A game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13744_ _07609_ _07610_ _07617_ net278 net241 vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__a221o_1
XANTENNA__10807__A2 _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17196__A1 _02387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10956_ game.CPU.applesa.ab.absxs.body_x\[117\] net321 vssd1 vssd1 vccd1 vccd1 _04846_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_63_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_317_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16463_ net214 _02417_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__nor2_4
X_19251_ clknet_leaf_7_clk _00065_ _00889_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11523__B net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13675_ game.writer.tracker.frame\[495\] net709 net672 game.writer.tracker.frame\[496\]
+ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__o22a_1
XANTENNA__16943__A1 _02379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10887_ net1172 net422 net417 net1170 _04788_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__o221a_1
XFILLER_0_195_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15414_ game.writer.updater.commands.count\[8\] game.writer.updater.commands.count\[7\]
+ _01441_ game.writer.updater.commands.count\[9\] game.writer.updater.commands.count\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__o311a_1
X_18202_ net580 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__inv_2
X_12626_ _06370_ _06371_ _06501_ _06502_ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__or4_2
X_19182_ clknet_leaf_5_clk _01301_ _00844_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_16394_ _02251_ _02307_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_193_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11768__B1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18133_ net583 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15345_ game.writer.updater.commands.count\[4\] game.writer.updater.commands.count\[3\]
+ _08886_ vssd1 vssd1 vccd1 vccd1 _08887_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_310_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12557_ game.CPU.applesa.ab.absxs.body_y\[85\] net523 net370 game.CPU.applesa.ab.absxs.body_x\[86\]
+ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13509__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15011__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19554__RESET_B net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18064_ net607 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__inv_2
X_11508_ game.CPU.applesa.ab.check_walls.above.walls\[2\] net768 vssd1 vssd1 vccd1
+ vccd1 _05397_ sky130_fd_sc_hd__xor2_2
XFILLER_0_312_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15276_ _08828_ _08829_ vssd1 vssd1 vccd1 vccd1 _08830_ sky130_fd_sc_hd__nand2_1
X_12488_ game.CPU.applesa.ab.absxs.body_x\[83\] net528 vssd1 vssd1 vccd1 vccd1 _06365_
+ sky130_fd_sc_hd__and2_1
XANTENNA__16171__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold108 game.writer.tracker.frame\[244\] vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_232_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12354__B net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17015_ _02507_ net89 _02675_ net1506 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[350\]
+ sky130_fd_sc_hd__a22o_1
Xhold119 game.writer.tracker.frame\[298\] vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14227_ game.CPU.applesa.ab.absxs.body_x\[43\] net1047 vssd1 vssd1 vccd1 vccd1 _08101_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_297_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11439_ _05317_ _05318_ _05327_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_74_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14158_ net1103 net883 _08030_ _08031_ net1 vssd1 vssd1 vccd1 vccd1 _08032_ sky130_fd_sc_hd__o221a_1
XANTENNA__17120__A1 _02369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10743__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_256_Right_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13109_ net284 _06955_ _06963_ _06971_ net241 vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__o221a_1
XANTENNA__13368__S0 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12370__A game.CPU.applesa.ab.absxs.body_x\[115\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18966_ net1199 _00110_ _00637_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_14089_ net956 game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1 vccd1
+ vccd1 _07963_ sky130_fd_sc_hd__xor2_1
XFILLER_0_253_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19535__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17917_ net590 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_146_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13693__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_321_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18897_ clknet_leaf_2_clk _00002_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_280_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1170 game.CPU.applesa.ab.YMAX\[2\] vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09361__A1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1181 net1182 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__buf_1
XANTENNA__09361__B2 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17848_ _08936_ _01430_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__or2_1
Xfanout1192 game.CPU.walls.rand_wall.good_spot vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16496__B _02441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16631__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_169_Left_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19685__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17779_ _03127_ _03129_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19303__D _00015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19518_ clknet_leaf_28_clk game.writer.tracker.next_frame\[113\] net1287 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[113\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_88_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_293_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19449_ clknet_leaf_48_clk game.writer.tracker.next_frame\[44\] net1294 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[44\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_347_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16934__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11471__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_307_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09202_ game.CPU.applesa.ab.check_walls.above.walls\[135\] vssd1 vssd1 vccd1 vccd1
+ _03451_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10049__B net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_335_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_332_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_307_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09133_ game.CPU.applesa.ab.check_walls.above.walls\[8\] vssd1 vssd1 vccd1 vccd1
+ _03382_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12420__A1 game.CPU.applesa.ab.absxs.body_y\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_322_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_301_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout318_A _05213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_178_Left_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09064_ game.CPU.applesa.ab.absxs.body_y\[36\] vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19065__CLK net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold620 game.writer.tracker.frame\[127\] vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout106_X net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold631 game.writer.tracker.frame\[22\] vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16304__X _02303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold642 game.writer.tracker.frame\[225\] vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13381__C1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold653 game.CPU.kyle.L1.cnt_20ms\[13\] vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 game.writer.tracker.frame\[505\] vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_246_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10734__A1 game.CPU.applesa.ab.absxs.body_y\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10734__B2 game.CPU.applesa.ab.absxs.body_y\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout687_A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_223_Right_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12280__A _06059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ net1130 net850 _04195_ vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__a21o_1
XANTENNA__14476__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16870__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09897_ _03812_ _03815_ _03970_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout854_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_187_Left_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09352__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18902__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09352__B2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15591__A game.CPU.applesa.ab.check_walls.above.walls\[34\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18675__Q game.CPU.applesa.ab.absxs.body_x\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10810_ game.CPU.applesa.ab.absxs.body_y\[119\] _04702_ vssd1 vssd1 vccd1 vccd1 _04729_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_16_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13987__A1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11790_ net824 net395 _05675_ _05258_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__o211a_1
XANTENNA__13987__B2 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_257_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12439__B net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10741_ net932 game.CPU.applesa.ab.absxs.body_y\[103\] net234 _04715_ vssd1 vssd1
+ vccd1 vccd1 _01042_ sky130_fd_sc_hd__a31o_1
XANTENNA__14494__X _08368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout907_X net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_270_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16853__C net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13460_ net515 _07327_ _07329_ net216 vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__a211o_1
XFILLER_0_192_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10672_ _03285_ net233 vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_326_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12726__Y _06600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12411_ game.CPU.applesa.ab.absxs.body_y\[55\] net365 net379 game.CPU.applesa.ab.absxs.body_x\[53\]
+ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_196_Left_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_358_Right_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_353_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_326_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19408__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ _06869_ _06871_ _07104_ _06884_ net507 net679 vssd1 vssd1 vccd1 vccd1 _07265_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_279_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12411__B2 game.CPU.applesa.ab.absxs.body_x\[53\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_152_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_211_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15130_ net1209 net1234 game.CPU.applesa.ab.check_walls.above.walls\[158\] vssd1
+ vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__and3_1
X_12342_ _03313_ net362 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16153__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17350__A1 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_287_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14164__A1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_346_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13598__S0 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15061_ net1217 net1244 game.CPU.applesa.ab.check_walls.above.walls\[89\] vssd1 vssd1
+ vccd1 vccd1 _00284_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12273_ _06051_ _06158_ _06053_ _06052_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__or4bb_1
XANTENNA__12175__B1 _06059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19558__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14012_ net940 net781 vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__nand2_1
XANTENNA__13911__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09764__A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ game.CPU.applesa.ab.absxs.body_y\[38\] net538 vssd1 vssd1 vccd1 vccd1 _05114_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_268_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13911__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10725__B2 game.CPU.applesa.ab.absxs.body_y\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18820_ clknet_leaf_2_clk _01211_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dfxtp_1
XANTENNA__09591__A1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_281_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11155_ game.CPU.applesa.ab.absxs.body_x\[51\] net407 vssd1 vssd1 vccd1 vccd1 _05045_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_235_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14467__A2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15664__A1 game.CPU.applesa.ab.check_walls.above.walls\[51\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16861__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ game.CPU.applesa.twoapples.start_enable game.CPU.applesa.enable_in game.CPU.applesa.twoapples.y_final\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__and3_1
XANTENNA__15664__B2 game.CPU.applesa.ab.check_walls.above.walls\[55\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_297_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18751_ clknet_leaf_59_clk _01168_ _00488_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[37\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11518__B net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15963_ _01968_ _01969_ _01970_ _01973_ vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__or4_1
X_11086_ game.CPU.applesa.ab.absxs.body_y\[62\] net401 vssd1 vssd1 vccd1 vccd1 _04976_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__16597__A game.writer.tracker.frame\[97\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13675__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18582__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17702_ game.CPU.walls.rand_wall.input2 _03522_ _03080_ net1206 vssd1 vssd1 vccd1
+ vccd1 _01307_ sky130_fd_sc_hd__o211a_1
XFILLER_0_262_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10037_ net1174 _03491_ _04243_ _04244_ _04224_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__a221o_1
X_14914_ net1174 _03489_ _08689_ _08690_ _08421_ vssd1 vssd1 vccd1 vccd1 _08691_ sky130_fd_sc_hd__a221o_1
XANTENNA__09343__B2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15894_ game.CPU.applesa.ab.absxs.body_y\[41\] net448 vssd1 vssd1 vccd1 vccd1 _01906_
+ sky130_fd_sc_hd__xnor2_1
X_18682_ clknet_leaf_8_clk _01099_ _00419_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_108_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14219__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_357_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17633_ net1421 _03035_ _03036_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__a21oi_1
XANTENNA__18585__Q game.CPU.applesa.ab.absxs.body_y\[50\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14845_ _08641_ _08642_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[6\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13225__S net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13978__A1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15006__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17169__A1 _02465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14776_ _08582_ _08584_ _08596_ vssd1 vssd1 vccd1 vccd1 _08597_ sky130_fd_sc_hd__or3b_1
X_17564_ net428 _02829_ _04256_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13978__B2 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11988_ net783 net296 net290 game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1
+ vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_141_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09456__A1_N net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11989__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19303_ clknet_leaf_65_clk _00015_ _00918_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.impossible
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13727_ game.writer.tracker.frame\[253\] game.writer.tracker.frame\[255\] game.writer.tracker.frame\[256\]
+ game.writer.tracker.frame\[254\] net981 net1032 vssd1 vssd1 vccd1 vccd1 _07601_
+ sky130_fd_sc_hd__mux4_1
X_16515_ net157 _02345_ _02456_ net727 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__o31a_1
XFILLER_0_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10939_ _04822_ _04823_ _04824_ _04825_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__a22o_1
XANTENNA__11453__A2 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16916__A1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17495_ game.CPU.walls.enable_in2 game.CPU.modea.Qa\[0\] vssd1 vssd1 vccd1 vccd1
+ _02924_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19234_ clknet_leaf_57_clk net1420 _00872_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.normal1.number\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16446_ net134 _02243_ _02405_ net734 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__o31a_1
X_13658_ game.writer.tracker.frame\[45\] game.writer.tracker.frame\[47\] game.writer.tracker.frame\[48\]
+ game.writer.tracker.frame\[46\] net970 net1002 vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12938__C1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12609_ _03301_ net369 net519 game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1
+ vccd1 vccd1 _06486_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_325_Right_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16377_ game.writer.tracker.frame\[32\] net734 _02352_ _02355_ vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[32\] sky130_fd_sc_hd__a31o_1
X_19165_ clknet_leaf_67_clk _01285_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count_luck\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13589_ net222 _07457_ _07462_ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18116_ net584 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__inv_2
X_15328_ game.CPU.applesa.twomode.number\[2\] _08866_ net757 vssd1 vssd1 vccd1 vccd1
+ _08872_ sky130_fd_sc_hd__a21o_1
X_19096_ net1178 _00134_ _00767_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[141\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16144__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12084__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18047_ net660 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__inv_2
X_15259_ game.CPU.kyle.L1.nextState\[2\] _08809_ _08810_ net2008 vssd1 vssd1 vccd1
+ vccd1 _08817_ sky130_fd_sc_hd__a22oi_4
XPHY_EDGE_ROW_200_Left_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09674__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13902__A1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13902__B2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13908__B game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__B2 game.CPU.applesa.ab.absxs.body_y\[50\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18925__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ _04054_ _04055_ _04061_ _04062_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__a211o_1
Xfanout407 net408 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_2
XFILLER_0_277_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout418 net420 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_4
XANTENNA__17891__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10613__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19998_ clknet_leaf_44_clk _01422_ net1299 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout429 _00293_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_2
XANTENNA__16852__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_253_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09751_ net912 game.CPU.applesa.ab.check_walls.above.walls\[24\] _03392_ net1094
+ _03993_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__a221o_1
XANTENNA__12469__A1 game.CPU.applesa.ab.absxs.body_x\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18949_ clknet_leaf_68_clk net1410 _00620_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11428__B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13666__B1 _07420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12469__B2 game.CPU.applesa.ab.absxs.body_y\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09682_ net1139 _03293_ _03294_ net1148 _03919_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__a221o_1
XANTENNA__16300__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11692__A2 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13135__S net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_334_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12259__B net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16907__A1 _02479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout435_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10652__B1 _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout58 net59 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_2
Xfanout69 _02331_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__buf_4
XFILLER_0_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_312_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout223_X net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1344_A net1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09116_ game.CPU.right_button.eD1.Q2 vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__inv_2
XANTENNA__19700__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10507__B _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09047_ game.CPU.applesa.ab.absxs.body_y\[94\] vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__inv_2
XANTENNA__15586__A game.CPU.applesa.ab.check_walls.above.walls\[32\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14490__A _08092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1132_X net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09584__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold450 game.writer.tracker.frame\[287\] vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 game.writer.tracker.frame\[411\] vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout971_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold472 game.writer.tracker.frame\[312\] vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12722__B _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11904__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17096__B1 _02700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold483 game.writer.tracker.frame\[102\] vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 game.writer.tracker.frame\[525\] vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout83_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13106__C1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_284_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout930 net931 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__buf_2
XFILLER_0_337_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout941 game.CPU.applesa.y\[3\] vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_4
XANTENNA__11338__B net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ net1120 net1121 _04172_ net1118 vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__a31o_1
Xfanout952 net957 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__buf_2
Xfanout963 net982 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_8
XANTENNA__14489__X _08363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_69_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout974 net976 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_4
XANTENNA__09325__A1 net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout985 net987 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09325__B2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12960_ _06780_ _06781_ net685 vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__mux2_1
XANTENNA__17306__A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_231_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_273_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11911_ net807 net393 net308 net806 _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__a221o_1
X_12891_ game.writer.tracker.frame\[58\] game.writer.tracker.frame\[59\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_231_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14630_ _08475_ _08476_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[15\]
+ sky130_fd_sc_hd__nor2_1
X_11842_ net790 net390 _05723_ _05724_ _05729_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14082__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_346_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14561_ net447 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.abduyd.next_wall\[5\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__11073__B net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12884__S net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ net571 _05459_ _05462_ _05660_ _05458_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__o2111a_1
XANTENNA__12737__X _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16209__X _02221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12632__B2 game.CPU.applesa.ab.absxs.body_y\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16300_ net214 net197 _02297_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__and3_4
X_13512_ net186 _07379_ _07380_ _07385_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__a22o_1
XANTENNA__17020__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17280_ net162 net114 _02343_ net735 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__o31a_1
XANTENNA__09759__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10724_ game.CPU.applesa.ab.absxs.body_y\[38\] _04642_ _04643_ game.CPU.applesa.ab.absxs.body_y\[34\]
+ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__a22o_1
X_14492_ _08299_ _08300_ _08152_ vssd1 vssd1 vccd1 vccd1 _08366_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16231_ net173 _02230_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__nor2_1
XFILLER_0_222_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_22_clk_X clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13443_ net701 _06931_ _07316_ net508 vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_299_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_190_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10655_ game.CPU.applesa.ab.absxs.body_x\[35\] _04696_ _04697_ game.CPU.applesa.ab.absxs.body_x\[31\]
+ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__a22o_1
XANTENNA__09478__B game.CPU.applesa.ab.check_walls.above.walls\[176\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14385__B2 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15582__B1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17976__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12185__A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11199__A1 game.CPU.applesa.ab.absxs.body_x\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_180_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11199__B2 game.CPU.applesa.ab.absxs.body_y\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16162_ _02073_ _02075_ _02076_ _02173_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__or4_1
XANTENNA__19380__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13374_ net492 _06710_ _07247_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__a21o_1
XANTENNA__17695__B net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload17 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_8
XANTENNA__16126__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload28 clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__clkinv_8
X_10586_ net1123 _04656_ _04594_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__o21ai_4
Xclkload39 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__inv_6
X_15113_ net1207 net1230 game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1
+ vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__and3_1
XANTENNA__14137__A1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12325_ _04210_ _04258_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__or2_4
XANTENNA__18948__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16093_ game.CPU.applesa.ab.absxs.body_y\[109\] net337 vssd1 vssd1 vccd1 vccd1 _02105_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__14137__B2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13345__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_clk_X clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19921_ clknet_leaf_33_clk game.writer.tracker.next_frame\[516\] net1302 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[516\] sky130_fd_sc_hd__dfrtp_1
X_15044_ net1219 net1244 game.CPU.applesa.ab.check_walls.above.walls\[72\] vssd1 vssd1
+ vccd1 vccd1 _00266_ sky130_fd_sc_hd__and3_1
X_12256_ _06045_ _06141_ _06043_ _06044_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__or4bb_1
XANTENNA__13896__B1 game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16104__B net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11207_ _03230_ net323 vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__xnor2_1
X_19852_ clknet_leaf_36_clk game.writer.tracker.next_frame\[447\] net1356 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[447\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_282_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12187_ net795 net547 vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__and2_1
XFILLER_0_207_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18803_ clknet_leaf_1_clk game.CPU.clock1.next_counter\[6\] _00540_ vssd1 vssd1 vccd1
+ vccd1 game.CPU.clock1.counter\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_247_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11138_ game.CPU.applesa.ab.absxs.body_y\[71\] net399 vssd1 vssd1 vccd1 vccd1 _05028_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__11248__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19783_ clknet_leaf_24_clk game.writer.tracker.next_frame\[378\] net1347 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[378\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15943__B net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_305_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16995_ _02455_ net120 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__nand2_4
XFILLER_0_207_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18734_ clknet_leaf_16_clk _01151_ _00471_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[104\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_143_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_250_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11069_ _04950_ _04951_ _04955_ _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__or4_1
X_15946_ _03401_ net270 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_0_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_250_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18665_ clknet_leaf_64_clk _01082_ _00402_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[87\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_203_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19204__Q game.CPU.applesa.ab.XMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15877_ _01883_ _01884_ _01886_ _01887_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__or4_1
XFILLER_0_188_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17616_ game.CPU.kyle.L1.cnt_20ms\[10\] _03023_ game.CPU.kyle.L1.cnt_20ms\[11\] vssd1
+ vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14828_ game.CPU.randy.f1.c1.count\[0\] game.CPU.randy.f1.c1.count\[1\] _04340_ vssd1
+ vssd1 vccd1 vccd1 _08631_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18596_ clknet_leaf_60_clk _01016_ _00333_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[73\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12079__B net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_230_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17547_ net1264 game.CPU.clock1.game_state\[0\] _02822_ vssd1 vssd1 vccd1 vccd1 _02973_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_82_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14759_ net54 _08579_ _08580_ vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_290_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_322_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09669__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19723__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17478_ _02884_ _02893_ _02896_ _02906_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__a31o_1
XANTENNA__17562__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19217_ net1167 _00019_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.normal1.counter
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16429_ net195 _02392_ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__nor2_2
XANTENNA__17886__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_332_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_305_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19148_ net1187 _00191_ _00819_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[193\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10937__A1 game.CPU.applesa.ab.absxs.body_x\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10937__B2 game.CPU.applesa.ab.absxs.body_y\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14128__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14128__B2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13919__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19873__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19079_ net1185 _00115_ _00750_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[124\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_93_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16014__B net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17078__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout204 net208 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout215 net217 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_243_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18510__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout226 net227 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_285_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11362__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout237 _02250_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_238_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09803_ net1147 game.CPU.applesa.ab.check_walls.above.walls\[109\] vssd1 vssd1 vccd1
+ vccd1 _04046_ sky130_fd_sc_hd__xor2_1
XANTENNA__11362__B2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout248 _06618_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_2
XANTENNA__15853__B _08429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11158__B net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout259 _05195_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_2
XFILLER_0_157_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_165_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09307__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16668__C _02434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_241_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09307__B2 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ net1146 _03346_ game.CPU.applesa.ab.absxs.body_y\[32\] net896 _03971_ vssd1
+ vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__a221o_1
XANTENNA__09851__B game.CPU.applesa.ab.absxs.body_x\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_213_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10997__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14469__B net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09665_ net1139 game.CPU.applesa.ab.absxs.body_y\[38\] vssd1 vssd1 vccd1 vccd1 _03908_
+ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout552_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A3 _04594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout173_X net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19114__Q game.CPU.applesa.ab.check_walls.above.walls\[159\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09596_ net1139 game.CPU.applesa.ab.absxs.body_y\[74\] vssd1 vssd1 vccd1 vccd1 _03839_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_328_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15800__B2 game.CPU.applesa.ab.absxs.body_x\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1082_X net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_254_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16210__D1 _01597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17796__A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11621__B net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09298__B game.CPU.applesa.ab.check_walls.above.walls\[81\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12378__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10440_ net1444 net848 _04168_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__a21o_1
XANTENNA__17305__A1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16108__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_249_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09794__A1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16659__A3 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ net1895 net850 _04200_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__a21o_1
XANTENNA__09794__B2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_343_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12110_ _05367_ _05996_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__or2_1
X_13090_ game.writer.tracker.frame\[234\] game.writer.tracker.frame\[235\] net1000
+ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout974_X net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12452__B net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_265_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13342__A2 _06654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12041_ net800 net295 _05926_ _05927_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__a211o_1
Xhold280 game.writer.tracker.frame\[254\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_291_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold291 game.writer.tracker.frame\[195\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10253__A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout86_X net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_207_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16816__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_284_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15763__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 net761 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout771 net772 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_8
X_15800_ game.CPU.applesa.ab.absxs.body_y\[51\] net433 net462 game.CPU.applesa.ab.absxs.body_x\[51\]
+ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__o2bb2a_1
Xfanout782 game.CPU.applesa.ab.check_walls.above.walls\[188\] vssd1 vssd1 vccd1 vccd1
+ net782 sky130_fd_sc_hd__buf_2
X_16780_ net152 _02452_ net107 _02595_ net1676 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[195\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_244_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13992_ net984 game.CPU.applesa.ab.check_walls.above.walls\[76\] vssd1 vssd1 vccd1
+ vccd1 _07866_ sky130_fd_sc_hd__xor2_1
Xfanout793 game.CPU.applesa.ab.check_walls.above.walls\[132\] vssd1 vssd1 vccd1 vccd1
+ net793 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14379__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12943_ net480 _06816_ _06815_ net223 vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__o211a_1
X_15731_ game.CPU.applesa.ab.absxs.body_x\[14\] net467 vssd1 vssd1 vccd1 vccd1 _01743_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16044__A1 game.CPU.applesa.ab.absxs.body_x\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16044__B2 game.CPU.applesa.ab.absxs.body_y\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_354_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ net652 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12874_ game.writer.tracker.frame\[8\] game.writer.tracker.frame\[9\] net1003 vssd1
+ vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__mux2_1
X_15662_ _03408_ net345 net443 net819 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__a22o_1
XANTENNA__19746__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18620__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12097__A2_N net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17401_ game.CPU.kyle.L1.nextState\[5\] game.CPU.kyle.L1.nextState\[4\] _02817_ vssd1
+ vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_202_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ game.CPU.clock1.counter\[9\] _08464_ net267 vssd1 vssd1 vccd1 vccd1 _08466_
+ sky130_fd_sc_hd__o21ai_1
X_11825_ game.CPU.applesa.ab.check_walls.above.walls\[124\] net390 vssd1 vssd1 vccd1
+ vccd1 _05713_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_276_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18381_ net596 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__inv_2
X_15593_ _03399_ game.CPU.walls.rand_wall.abduyd.next_wall\[4\] net433 game.CPU.applesa.ab.check_walls.above.walls\[39\]
+ _01604_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__a221o_1
XFILLER_0_358_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13802__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17332_ game.writer.updater.commands.mode\[1\] _01579_ net576 vssd1 vssd1 vccd1 vccd1
+ _02765_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_218_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _08413_ _08415_ _04257_ vssd1 vssd1 vccd1 vccd1 _08416_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09489__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11756_ game.CPU.applesa.ab.check_walls.above.walls\[174\] net300 _05637_ _05643_
+ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_327_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10707_ _03337_ net425 vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__nor2_1
X_17263_ net207 net112 _02393_ _02746_ net1604 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[527\]
+ sky130_fd_sc_hd__a32o_1
X_14475_ _03292_ net1074 net1056 _03290_ vssd1 vssd1 vccd1 vccd1 _08349_ sky130_fd_sc_hd__o22a_1
XANTENNA__18770__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15003__B net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19896__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11687_ net744 _05568_ _05569_ net567 _05575_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19002_ net1189 _00229_ _00673_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_299_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13426_ _07298_ _07299_ net477 vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__mux2_1
XANTENNA__09776__X _04019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16214_ _02163_ _02172_ _02175_ _02225_ vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__nand4_1
X_17194_ _02502_ net75 _02729_ net1566 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[475\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10638_ net1269 _04630_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_314_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19694__Q game.writer.tracker.frame\[289\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_342_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16145_ _03438_ net451 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__xnor2_1
X_13357_ _06665_ _06675_ net688 vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__mux2_1
XANTENNA__09936__B net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10569_ _04591_ _04617_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__nand2_2
XFILLER_0_140_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13318__C1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19126__CLK net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_307_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12308_ _06027_ _06193_ _06029_ _06028_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__or4bb_1
X_16076_ game.CPU.applesa.ab.absxs.body_y\[86\] net438 vssd1 vssd1 vccd1 vccd1 _02088_
+ sky130_fd_sc_hd__xnor2_1
X_13288_ net186 _07072_ _07103_ _07161_ net178 vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_287_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12362__B net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13869__B1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19904_ clknet_leaf_20_clk game.writer.tracker.next_frame\[499\] net1316 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[499\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_267_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15027_ net1222 net1250 net818 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__and3_1
XANTENNA__15954__A game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12239_ game.CPU.applesa.ab.check_walls.above.walls\[150\] net417 vssd1 vssd1 vccd1
+ vccd1 _06125_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09537__B2 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_229_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10163__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18330__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12541__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15592__A2_N game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19835_ clknet_leaf_33_clk game.writer.tracker.next_frame\[430\] net1325 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[430\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_208_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15673__B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19276__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13474__A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17267__A1_N net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_272_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13097__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16822__A3 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19766_ clknet_leaf_29_clk game.writer.tracker.next_frame\[361\] net1291 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[361\] sky130_fd_sc_hd__dfrtp_1
X_16978_ _02252_ net167 _02664_ net717 vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__o31a_2
XANTENNA__14294__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 gpio_in[2] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_18717_ clknet_leaf_66_clk _01134_ _00454_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[83\]
+ sky130_fd_sc_hd__dfrtp_4
X_15929_ net795 net444 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__xnor2_1
X_19697_ clknet_leaf_29_clk game.writer.tracker.next_frame\[292\] net1284 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[292\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17232__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09450_ _03686_ _03688_ _03691_ _03692_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__and4_1
X_18648_ clknet_leaf_12_clk _01065_ _00385_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[54\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_318_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18773__Q game.CPU.applesa.ab.absxs.body_x\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09381_ net1112 _03382_ _03384_ net1160 vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__a22o_1
X_18579_ clknet_leaf_53_clk _00999_ _00316_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[40\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15794__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09399__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload72_A clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16009__B net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12537__B net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16889__A3 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13021__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13021__B2 _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09776__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09776__B2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout300_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_329_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12272__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19619__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15864__A game.CPU.applesa.ab.absxs.body_y\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11169__A game.CPU.applesa.ab.absxs.body_y\[76\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18240__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1307_A net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16679__B _02237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12532__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09862__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout767_A game.CPU.applesa.ab.apple_possible\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19769__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14285__B1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18643__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14199__B net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ net1125 game.CPU.applesa.ab.absxs.body_y\[87\] vssd1 vssd1 vccd1 vccd1 _03960_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__13183__S1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11616__B net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_260_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout934_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09700__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__B2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ _03887_ _03888_ _03889_ _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__or4b_1
XANTENNA__16577__A2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_334_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14588__B2 net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12287__X _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ net922 game.CPU.applesa.ab.check_walls.above.walls\[42\] game.CPU.applesa.ab.check_walls.above.walls\[46\]
+ net904 vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__o22a_1
XANTENNA__18793__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12599__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11632__A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ net804 net316 net253 game.CPU.applesa.ab.check_walls.above.walls\[100\] vssd1
+ vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12590_ game.CPU.applesa.ab.absxs.body_x\[90\] net370 net359 game.CPU.applesa.ab.absxs.body_y\[88\]
+ _06324_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__a221o_1
XFILLER_0_355_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12447__B net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09102__A game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11541_ game.CPU.applesa.ab.check_walls.above.walls\[145\] net769 vssd1 vssd1 vccd1
+ vccd1 _05430_ sky130_fd_sc_hd__xor2_1
XANTENNA__11351__B net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10248__A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11810__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ net1267 net890 net987 _03302_ vssd1 vssd1 vccd1 vccd1 _08134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_279_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11472_ net828 net256 _05348_ _05360_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__o211a_1
XFILLER_0_269_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08941__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15758__B net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13211_ net704 _07084_ _07081_ net230 vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__o211a_1
X_10423_ game.CPU.right_button.eD1.Q1 _03365_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__nand2_1
XANTENNA__09767__A1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_213_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14191_ game.CPU.applesa.ab.absxs.body_y\[96\] net1042 vssd1 vssd1 vccd1 vccd1 _08065_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__09767__B2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ game.writer.tracker.frame\[152\] game.writer.tracker.frame\[153\] net1035
+ vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_249_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10354_ game.CPU.walls.rand_wall.counter2\[4\] _04516_ _04519_ vssd1 vssd1 vccd1
+ vccd1 _04520_ sky130_fd_sc_hd__a21boi_1
XANTENNA__19299__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12182__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19019__Q game.CPU.applesa.ab.check_walls.above.walls\[64\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_295_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13073_ _06943_ _06944_ _06946_ _06945_ net491 net687 vssd1 vssd1 vccd1 vccd1 _06947_
+ sky130_fd_sc_hd__mux4_2
X_17950_ net614 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__inv_2
X_10285_ _03214_ net1436 _04473_ _04475_ vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__o31a_1
X_16901_ _02237_ _02272_ _02311_ net556 vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a31oi_2
XTAP_TAPCELL_ROW_111_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12024_ game.CPU.applesa.ab.check_walls.above.walls\[14\] net290 vssd1 vssd1 vccd1
+ vccd1 _05911_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15493__B _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17881_ net656 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_228_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19620_ clknet_leaf_23_clk game.writer.tracker.next_frame\[215\] net1337 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[215\] sky130_fd_sc_hd__dfrtp_1
X_16832_ net145 _02369_ net102 _02610_ net1488 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[230\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__16804__A3 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_302_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14276__B1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_272_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout590 net591 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__buf_4
XFILLER_0_217_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19551_ clknet_leaf_34_clk game.writer.tracker.next_frame\[146\] net1328 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[146\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_205_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16763_ net168 _02331_ net65 _02590_ net1740 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[183\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_205_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_224_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13975_ net949 game.CPU.applesa.ab.check_walls.above.walls\[86\] vssd1 vssd1 vccd1
+ vccd1 _07849_ sky130_fd_sc_hd__or2_1
X_18502_ net601 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__inv_2
XFILLER_0_244_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_232_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload9_A clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15714_ game.CPU.applesa.ab.absxs.body_y\[11\] net435 vssd1 vssd1 vccd1 vccd1 _01726_
+ sky130_fd_sc_hd__xnor2_1
X_19482_ clknet_leaf_18_clk game.writer.tracker.next_frame\[77\] net1308 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[77\] sky130_fd_sc_hd__dfrtp_1
X_12926_ net220 _06797_ _06799_ net282 vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__a31o_1
X_16694_ net204 net53 net61 _02564_ net1452 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[140\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_319_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_244_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18433_ net586 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__inv_2
XFILLER_0_347_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15776__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15645_ game.CPU.applesa.ab.check_walls.above.walls\[74\] net466 vssd1 vssd1 vccd1
+ vccd1 _01657_ sky130_fd_sc_hd__xnor2_1
X_12857_ game.writer.tracker.frame\[302\] game.writer.tracker.frame\[303\] net989
+ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11542__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15014__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18364_ net596 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ net817 net393 net302 game.CPU.applesa.ab.check_walls.above.walls\[62\] _05695_
+ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__a221o_1
X_12788_ game.writer.tracker.frame\[380\] game.writer.tracker.frame\[381\] net1034
+ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15576_ _03429_ net339 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_196_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12357__B net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10065__A1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17315_ net1768 _02761_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[564\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__15528__A0 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14527_ _08399_ _08400_ _07742_ vssd1 vssd1 vccd1 vccd1 _08401_ sky130_fd_sc_hd__a21bo_1
X_11739_ game.CPU.applesa.ab.check_walls.above.walls\[157\] net305 vssd1 vssd1 vccd1
+ vccd1 _05627_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18295_ net641 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_313_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17019__A2_N net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18325__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17246_ _02275_ _02448_ _02742_ net1731 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[514\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14458_ game.CPU.applesa.ab.absxs.body_x\[14\] net1056 vssd1 vssd1 vccd1 vccd1 _08332_
+ sky130_fd_sc_hd__or2_1
XANTENNA__15668__B net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13409_ _06873_ _06887_ net680 vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__mux2_1
X_17177_ _02475_ net73 _02725_ net1825 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[462\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14389_ game.CPU.applesa.ab.absxs.body_x\[4\] net890 net884 game.CPU.applesa.ab.absxs.body_x\[5\]
+ _08259_ vssd1 vssd1 vccd1 vccd1 _08263_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16128_ game.CPU.applesa.ab.check_walls.above.walls\[160\] net354 net450 game.CPU.applesa.ab.check_walls.above.walls\[164\]
+ _01666_ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_77_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12092__B net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_269_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08950_ net1141 vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__inv_2
X_16059_ game.CPU.applesa.ab.check_walls.above.walls\[197\] net445 vssd1 vssd1 vccd1
+ vccd1 _02071_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_90_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18666__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12514__B1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19911__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17048__A3 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16256__A1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_324_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19818_ clknet_leaf_37_clk game.writer.tracker.next_frame\[413\] net1350 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[413\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_285_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19931__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10621__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10540__A2 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Left_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_263_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13165__S1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19749_ clknet_leaf_24_clk game.writer.tracker.next_frame\[344\] net1341 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[344\] sky130_fd_sc_hd__dfrtp_1
X_09502_ net916 game.CPU.applesa.ab.check_walls.above.walls\[49\] game.CPU.applesa.ab.check_walls.above.walls\[51\]
+ net926 _03744_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13490__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_338_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09433_ net927 game.CPU.applesa.ab.absxs.body_x\[59\] _03340_ net1160 vssd1 vssd1
+ vccd1 vccd1 _03676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15767__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout250_A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12548__A game.CPU.applesa.ab.absxs.body_y\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09364_ _03601_ _03602_ _03603_ _03605_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__or4_1
XFILLER_0_304_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12557__A2_N net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11171__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15519__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15859__A game.CPU.applesa.ab.absxs.body_x\[115\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_129_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_20 _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09295_ net1146 _03425_ _03426_ net1128 vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout515_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_31 _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout136_X net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_42 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09857__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16192__B1 _02200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15578__B net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16731__A2 _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_320_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19441__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11556__A1 _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_X net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__B2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout884_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_249_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1212_X net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_262_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19591__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17039__A3 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ _04276_ _04277_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_345_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19601__RESET_B net1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11346__B net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout937_X net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ game.writer.tracker.frame\[130\] net841 net834 game.writer.tracker.frame\[129\]
+ vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__o22a_1
XFILLER_0_214_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10972_ game.CPU.applesa.ab.absxs.body_y\[75\] net397 vssd1 vssd1 vccd1 vccd1 _04862_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_281_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap66 _02514_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_4
X_12711_ net1065 net1057 net1048 vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_356_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13691_ game.writer.tracker.frame\[510\] net843 net837 game.writer.tracker.frame\[509\]
+ vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__o22a_1
XFILLER_0_329_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17211__A3 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13053__S net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_273_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15430_ _01434_ _01432_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__nand2b_1
X_12642_ game.CPU.applesa.ab.absxs.body_x\[18\] net371 game.CPU.applesa.twoapples.absxs.next_head\[4\]
+ _03354_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__a22o_1
XFILLER_0_214_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16970__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__Y _04442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_215_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15361_ game.writer.updater.commands.cmd_num\[2\] _08877_ _08897_ _08902_ vssd1 vssd1
+ vccd1 vccd1 _08903_ sky130_fd_sc_hd__o22a_2
X_12573_ game.CPU.applesa.ab.absxs.body_y\[18\] net519 net360 game.CPU.applesa.ab.absxs.body_y\[16\]
+ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_343_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17100_ _02497_ net60 _02702_ net1987 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[408\]
+ sky130_fd_sc_hd__a22o_1
X_14312_ game.CPU.applesa.ab.absxs.body_y\[56\] net871 net859 game.CPU.applesa.ab.absxs.body_y\[59\]
+ _08185_ vssd1 vssd1 vccd1 vccd1 _08186_ sky130_fd_sc_hd__a221o_1
X_11524_ _05412_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__inv_2
X_18080_ net669 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__inv_2
X_15292_ game.CPU.applesa.twomode.number\[4\] game.CPU.applesa.twomode.counter_flip
+ vssd1 vssd1 vccd1 vccd1 _08842_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_324_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_237_Right_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_230_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17031_ _02375_ net85 _02681_ net1697 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[360\]
+ sky130_fd_sc_hd__a22o_1
X_14243_ _08114_ _08115_ _08116_ vssd1 vssd1 vccd1 vccd1 _08117_ sky130_fd_sc_hd__or3_2
X_11455_ game.CPU.applesa.ab.check_walls.above.walls\[76\] net253 net260 game.CPU.applesa.ab.check_walls.above.walls\[79\]
+ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12193__A game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10406_ _04341_ _04549_ _04552_ _04553_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__a211oi_1
X_14174_ _03252_ net1050 net858 game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1
+ vccd1 vccd1 _08048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17278__A3 _02341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11386_ game.CPU.applesa.ab.check_walls.above.walls\[181\] net318 _05270_ _05272_
+ _05274_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__o2111a_1
XANTENNA__15000__C net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13125_ _06997_ _06998_ net504 vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10337_ _04487_ _04510_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__nand2_1
X_18982_ net1201 _00207_ _00653_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_284_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14497__B1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10770__A2 _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13056_ game.writer.tracker.frame\[224\] game.writer.tracker.frame\[225\] net1011
+ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_226_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ net660 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__inv_2
X_10268_ _03493_ net746 vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__nand2_1
XANTENNA__16238__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16112__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1330 net1331 vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__clkbuf_4
X_12007_ _05891_ _05892_ _05893_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__or3_2
Xfanout1341 net1359 vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__clkbuf_2
XANTENNA__15009__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1352 net1353 vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_292_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17864_ _01443_ _03173_ _03184_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__o21bai_1
X_10199_ net1082 _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__and2_1
XANTENNA__16789__A2 _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19603_ clknet_leaf_19_clk game.writer.tracker.next_frame\[198\] net1342 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[198\] sky130_fd_sc_hd__dfrtp_1
X_16815_ _02506_ net105 _02604_ net1897 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[221\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_255_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09007__A game.CPU.applesa.ab.absxs.body_x\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17795_ _06556_ _03134_ _03136_ net721 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__a22o_1
XANTENNA__15997__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19534_ clknet_leaf_32_clk game.writer.tracker.next_frame\[129\] net1291 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[129\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_198_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16746_ net163 net53 net101 _02584_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[172\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13958_ net1054 game.CPU.applesa.ab.check_walls.above.walls\[178\] vssd1 vssd1 vccd1
+ vccd1 _07832_ sky130_fd_sc_hd__xor2_1
X_12909_ net510 _06666_ _06668_ net228 vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__o211a_1
X_19465_ clknet_leaf_40_clk game.writer.tracker.next_frame\[60\] net1358 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[60\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16677_ net1981 _02554_ _02555_ _02448_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[130\]
+ sky130_fd_sc_hd__a22o_1
X_13889_ net950 game.CPU.applesa.ab.check_walls.above.walls\[102\] vssd1 vssd1 vccd1
+ vccd1 _07763_ sky130_fd_sc_hd__or2_1
XANTENNA__12368__A game.CPU.applesa.ab.absxs.body_y\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18416_ net626 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
X_15628_ _03482_ net336 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_237_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19396_ clknet_leaf_55_clk net1386 net1280 vssd1 vssd1 vccd1 vccd1 game.writer.control.button5.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14421__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15679__A _03385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18347_ net594 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__inv_2
X_15559_ _08924_ _08927_ net576 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__or3_1
XANTENNA__10589__A2 _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12983__B1 _06856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ game.CPU.applesa.ab.absxs.body_y\[82\] vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09677__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18278_ net645 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_204_Right_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17229_ _02412_ net123 net121 _02738_ net1829 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[501\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_287_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17269__A3 _02486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_326_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload35_A clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13927__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09982_ game.CPU.applesa.off_bc.Q2 game.CPU.applesa.off_bc.Q1 vssd1 vssd1 vccd1 vccd1
+ _04208_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_228_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16303__A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10761__A2 _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12550__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16022__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout298_A _05858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11447__A game.CPU.applesa.ab.check_walls.above.walls\[73\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1005_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13138__S1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15861__B net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout465_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_337_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_339_Right_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20055__1373 vssd1 vssd1 vccd1 vccd1 _20055__1373/HI net1373 sky130_fd_sc_hd__conb_1
XFILLER_0_189_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12278__A net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout253_X net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19807__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09416_ net1091 game.CPU.applesa.ab.absxs.body_x\[98\] vssd1 vssd1 vccd1 vccd1 _03659_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_121_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14412__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16952__A2 _02638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18961__Q game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09347_ net1093 game.CPU.applesa.ab.absxs.body_x\[10\] vssd1 vssd1 vccd1 vccd1 _03590_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__13766__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_353_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09278_ game.CPU.applesa.normal1.counter_normal vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19957__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16704__A2 _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12725__B net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10526__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11240_ _03258_ net320 vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_210_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12821__S0 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout887_X net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ game.CPU.applesa.ab.absxs.body_x\[76\] net324 vssd1 vssd1 vccd1 vccd1 _05061_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_132_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14479__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16213__A _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10752__A2 _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10122_ net1166 net851 game.CPU.applesa.ab.good_collision _03214_ vssd1 vssd1 vccd1
+ vccd1 _01339_ sky130_fd_sc_hd__a211o_1
XANTENNA__12460__B net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__Y _04639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13151__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11357__A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ game.CPU.applesa.twoapples.count_luck\[1\] game.CPU.applesa.twoapples.count_luck\[0\]
+ game.CPU.applesa.twoapples.count_luck\[2\] vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__a21o_1
X_14930_ _08680_ _08683_ _08706_ _08664_ vssd1 vssd1 vccd1 vccd1 _08707_ sky130_fd_sc_hd__a211o_1
XFILLER_0_356_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_261_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19337__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10504__A2 _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11701__B2 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11076__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A2 game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12887__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15771__B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ game.CPU.randy.f1.c1.count\[13\] game.CPU.randy.f1.c1.count\[14\] _08649_
+ vssd1 vssd1 vccd1 vccd1 _08651_ sky130_fd_sc_hd__and3_1
X_16600_ _02345_ _02513_ _02511_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[97\]
+ sky130_fd_sc_hd__o21ai_1
X_13812_ game.writer.tracker.frame\[409\] game.writer.tracker.frame\[411\] game.writer.tracker.frame\[412\]
+ game.writer.tracker.frame\[410\] net980 net1035 vssd1 vssd1 vccd1 vccd1 _07686_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_221_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17580_ game.CPU.kyle.L1.cnt_20ms\[2\] game.CPU.kyle.L1.cnt_20ms\[1\] game.CPU.kyle.L1.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__and3_1
XFILLER_0_202_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14792_ game.CPU.randy.counter1.count\[4\] _08604_ game.CPU.randy.counter1.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _08609_ sky130_fd_sc_hd__a21o_1
XANTENNA__09658__B1 game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14387__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16531_ net146 net125 _02467_ _02463_ net1916 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[74\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_329_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13743_ _07613_ _07616_ net228 vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__mux2_1
XANTENNA__19487__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_306_Right_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10955_ _03286_ net319 vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11804__B net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19250_ clknet_leaf_7_clk _00064_ _00888_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13206__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16462_ net242 _02285_ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__or2_2
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13674_ _07546_ _07547_ net477 vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__mux2_1
XANTENNA__14403__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10886_ net1170 net417 net547 net1171 _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__a221o_1
XFILLER_0_344_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18201_ net580 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__inv_2
X_15413_ game.writer.updater.commands.count\[2\] _08887_ game.writer.updater.commands.count\[6\]
+ game.writer.updater.commands.count\[5\] vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__o211a_1
XFILLER_0_356_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13757__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12625_ _06363_ _06368_ _06369_ _06372_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__or4_1
X_19181_ clknet_leaf_5_clk _01300_ _00843_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_16393_ net1972 net720 _02366_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[37\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__12916__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_193_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11768__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18132_ net578 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__inv_2
XANTENNA__11768__B2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09497__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15344_ game.writer.updater.commands.count\[1\] game.writer.updater.commands.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08886_ sky130_fd_sc_hd__or2_1
X_12556_ game.CPU.applesa.ab.absxs.body_y\[86\] net517 net523 game.CPU.applesa.ab.absxs.body_y\[85\]
+ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_310_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ game.CPU.applesa.ab.check_walls.above.walls\[5\] net317 vssd1 vssd1 vccd1
+ vccd1 _05396_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_10_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18063_ net607 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__inv_2
XANTENNA__15011__B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12487_ game.CPU.applesa.ab.absxs.body_x\[83\] net528 vssd1 vssd1 vccd1 vccd1 _06364_
+ sky130_fd_sc_hd__nor2_1
X_15275_ _08816_ _08818_ vssd1 vssd1 vccd1 vccd1 _08829_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_232_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_297_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17014_ _02506_ net89 _02675_ net1848 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[349\]
+ sky130_fd_sc_hd__a22o_1
Xhold109 game.CPU.applesa.ab.apple_location\[5\] vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_312_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11438_ net568 _05319_ _05322_ net744 _05326_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__o221a_1
XFILLER_0_151_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14226_ game.CPU.applesa.ab.absxs.body_x\[43\] net1047 vssd1 vssd1 vccd1 vccd1 _08100_
+ sky130_fd_sc_hd__or2_1
XANTENNA__15946__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_297_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14157_ net1141 net955 vssd1 vssd1 vccd1 vccd1 _08031_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_74_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11369_ net777 _05257_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_238_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10743__A2 game.CPU.applesa.ab.absxs.body_y\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13108_ net280 _06980_ _06981_ net246 vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__o31a_1
X_18965_ net1200 _00099_ _00636_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_14088_ _07957_ _07958_ _07959_ _07961_ vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__nor4_1
XANTENNA__12370__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19207__Q game.CPU.applesa.ab.YMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13039_ net697 _06871_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__or2_1
XFILLER_0_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17916_ net605 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__inv_2
XFILLER_0_265_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_266_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18896_ clknet_leaf_2_clk _00001_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_146_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_321_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1160 net1161 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__clkbuf_8
Xfanout1171 game.CPU.applesa.ab.YMAX\[1\] vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__clkbuf_4
X_17847_ game.writer.updater.commands.count\[10\] _03169_ vssd1 vssd1 vccd1 vccd1
+ _03172_ sky130_fd_sc_hd__and2_1
Xfanout1182 net1183 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__clkbuf_2
XANTENNA__15681__B net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18704__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1193 net1194 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__buf_2
XANTENNA__16631__A1 _02237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17778_ game.CPU.applesa.twoapples.count\[2\] game.CPU.applesa.twoapples.count\[1\]
+ game.CPU.applesa.twoapples.count\[3\] _03127_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__nand4_2
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19517_ clknet_leaf_28_clk game.writer.tracker.next_frame\[112\] net1287 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[112\] sky130_fd_sc_hd__dfrtp_1
X_16729_ _02512_ net63 _02578_ game.writer.tracker.frame\[161\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[161\] sky130_fd_sc_hd__a22o_1
XFILLER_0_76_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11714__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17889__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17187__A2 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_347_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19448_ clknet_leaf_47_clk game.writer.tracker.next_frame\[43\] net1294 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[43\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18854__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16934__A2 _02524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09201_ game.CPU.applesa.ab.check_walls.above.walls\[134\] vssd1 vssd1 vccd1 vccd1
+ _03450_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19379_ net1165 _01385_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twomode.counter_flip
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_157_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_332_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09132_ net831 vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12420__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16698__A1 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14158__C1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09200__A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16017__B net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ game.CPU.applesa.ab.absxs.body_y\[37\] vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout213_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18513__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_303_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold610 game.writer.tracker.frame\[13\] vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold621 game.writer.tracker.frame\[57\] vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_288_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold632 game.writer.tracker.frame\[420\] vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 game.writer.tracker.frame\[387\] vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_330_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold654 game.writer.tracker.frame\[7\] vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 game.writer.tracker.frame\[551\] vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16033__A game.CPU.applesa.ab.absxs.body_x\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17111__A2 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1122_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_246_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09965_ net1128 _04193_ _04194_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_51_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16870__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__A game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_243_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09896_ _04113_ _04117_ _04138_ _03857_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__o211a_2
XANTENNA__09888__B1 _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_X net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10512__C net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18956__Q game.CPU.applesa.ab.check_walls.above.walls\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09352__A2 game.CPU.applesa.ab.absxs.body_x\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15591__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout468_X net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13392__A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16622__A1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_257_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ game.CPU.applesa.ab.absxs.body_y\[107\] _04658_ vssd1 vssd1 vccd1 vccd1 _04715_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_270_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18691__Q game.CPU.applesa.ab.absxs.body_x\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10671_ _04594_ _04656_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__nand2_2
XANTENNA__12736__A _06607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ game.CPU.applesa.ab.absxs.body_x\[53\] net379 net525 game.CPU.applesa.ab.absxs.body_y\[53\]
+ _06286_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_24_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13390_ _07260_ _07263_ net206 vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_313_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16689__A1 _02464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12341_ net359 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.absxs.next_head\[4\]
+ sky130_fd_sc_hd__inv_6
XANTENNA__17350__A2 _02779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15060_ net1217 net1246 game.CPU.applesa.ab.check_walls.above.walls\[88\] vssd1 vssd1
+ vccd1 vccd1 _00283_ sky130_fd_sc_hd__and3_1
XANTENNA__14164__A2 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12272_ game.CPU.applesa.ab.check_walls.above.walls\[157\] net548 vssd1 vssd1 vccd1
+ vccd1 _06158_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_287_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14011_ net948 game.CPU.applesa.ab.check_walls.above.walls\[190\] vssd1 vssd1 vccd1
+ vccd1 _07885_ sky130_fd_sc_hd__xor2_1
XANTENNA__16214__Y _00288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12175__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11223_ game.CPU.applesa.ab.absxs.body_y\[38\] net540 vssd1 vssd1 vccd1 vccd1 _05113_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_268_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_281_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11154_ _05032_ _05036_ _05040_ _05043_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__or4_4
XANTENNA__12190__B net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18727__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16861__A1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10105_ game.CPU.applesa.twoapples.start_enable game.CPU.applesa.enable_in vssd1
+ vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__nand2_1
XANTENNA__15664__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18750_ clknet_leaf_59_clk _01167_ _00487_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[36\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__15782__A game.CPU.applesa.ab.absxs.body_y\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_297_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11085_ _03238_ net406 vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__xnor2_1
X_15962_ _01964_ _01965_ _01971_ _01972_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__or4_1
XANTENNA__12478__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__B1 _04032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17701_ _03076_ _03077_ _03078_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__nand3_2
X_10036_ game.CPU.applesa.ab.XMAX\[1\] _04210_ _04232_ net1174 vssd1 vssd1 vccd1 vccd1
+ _04244_ sky130_fd_sc_hd__o22a_1
X_14913_ game.CPU.applesa.ab.XMAX\[1\] _08417_ _08419_ net1174 vssd1 vssd1 vccd1 vccd1
+ _08690_ sky130_fd_sc_hd__o22a_1
X_18681_ clknet_leaf_12_clk _01098_ _00418_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[119\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_236_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15893_ game.CPU.applesa.ab.absxs.body_x\[40\] net273 vssd1 vssd1 vccd1 vccd1 _01905_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_349_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17632_ net1421 _03035_ net429 vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__o21ai_1
X_14844_ game.CPU.randy.f1.c1.count\[6\] _08638_ vssd1 vssd1 vccd1 vccd1 _08642_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_357_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18877__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16884__Y _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17563_ _04484_ _02825_ _02833_ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__and3_1
XANTENNA__13978__A2 game.CPU.applesa.ab.check_walls.above.walls\[80\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15006__B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14775_ game.CPU.randy.counter1.count\[12\] game.CPU.randy.counter1.count\[8\] game.CPU.randy.counter1.count\[1\]
+ net265 vssd1 vssd1 vccd1 vccd1 _08596_ sky130_fd_sc_hd__a31o_1
XFILLER_0_175_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11987_ _05870_ _05871_ _05873_ _05869_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__a211o_1
X_19302_ clknet_leaf_56_clk game.CPU.applesa.ab.check_walls.above.collision _00917_
+ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.collision_up sky130_fd_sc_hd__dfrtp_1
X_16514_ net222 _02244_ net236 net195 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__or4_4
XFILLER_0_252_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13726_ net210 _07593_ _07599_ net277 vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__o211a_1
X_10938_ game.CPU.applesa.ab.absxs.body_x\[10\] net409 net398 game.CPU.applesa.ab.absxs.body_y\[11\]
+ _04821_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__o221a_1
X_17494_ game.CPU.walls.enable_in2 game.CPU.modea.Qa\[0\] vssd1 vssd1 vccd1 vccd1
+ _02923_ sky130_fd_sc_hd__nor2_1
XANTENNA__16916__A2 _02643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19233_ clknet_leaf_57_clk net1427 _00871_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.normal1.number\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16445_ _02321_ net166 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_234_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13657_ _07527_ _07530_ net205 vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__mux2_1
X_10869_ _04768_ _04769_ _04771_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__nor3_1
XFILLER_0_317_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12608_ _06379_ _06380_ _06482_ _06484_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__or4_1
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19164_ clknet_leaf_67_clk _01284_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count_luck\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_16376_ net137 _02258_ _02354_ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__and3_1
X_13588_ net213 _07461_ net283 vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__a21o_1
X_18115_ net584 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15957__A game.CPU.applesa.ab.check_walls.above.walls\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15327_ game.CPU.applesa.twomode.number\[2\] _08866_ vssd1 vssd1 vccd1 vccd1 _08871_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11610__B1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19095_ net1177 _00133_ _00766_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[140\]
+ sky130_fd_sc_hd__dfrtp_4
X_12539_ game.CPU.applesa.ab.absxs.body_x\[42\] net371 net526 game.CPU.applesa.ab.absxs.body_y\[41\]
+ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__o22ai_1
XANTENNA__12933__X _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19502__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18046_ net660 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19704__RESET_B net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15676__B net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15258_ game.CPU.kyle.L1.currentState\[0\] net1259 _08808_ vssd1 vssd1 vccd1 vccd1
+ _08816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_297_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14209_ game.CPU.applesa.ab.absxs.body_x\[95\] net1044 vssd1 vssd1 vccd1 vccd1 _08083_
+ sky130_fd_sc_hd__xor2_1
X_20054__1372 vssd1 vssd1 vccd1 vccd1 _20054__1372/HI net1372 sky130_fd_sc_hd__conb_1
XANTENNA__09674__B net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15189_ game.CPU.walls.enable_in2 _08761_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_285_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10716__A2 _04609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout408 game.CPU.applesa.ab.absxs.next_head\[3\] vssd1 vssd1 vccd1 vccd1 net408
+ sky130_fd_sc_hd__buf_4
X_19997_ clknet_leaf_44_clk _01421_ net1304 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[12\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout419 net420 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_4
XFILLER_0_277_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10613__B _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19652__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13764__X _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15692__A game.CPU.applesa.ab.absxs.body_x\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_265_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09750_ net1141 game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1 vccd1
+ vccd1 _03993_ sky130_fd_sc_hd__xor2_1
XANTENNA__13666__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_265_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12469__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18948_ clknet_leaf_68_clk net1405 _00619_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__15821__A2_N net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09690__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11677__B1 _05565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09681_ _03917_ _03918_ _03922_ _03923_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__a22o_1
X_18879_ clknet_leaf_5_clk game.CPU.randy.f1.c1.innerCount\[9\] _00574_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13416__S net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13418__A1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_240_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16122__A1_N game.CPU.applesa.ab.absxs.body_x\[54\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Left_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11444__B net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_334_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18508__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13940__A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout59 net60 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_2
XANTENNA__19400__Q game.CPU.applesa.x\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1072_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12929__B1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09578__A1_N net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11460__A game.CPU.applesa.ab.check_walls.above.walls\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_312_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12275__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09115_ game.writer.updater.commands.mode\[1\] vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16315__X _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13029__S0 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout216_X net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18243__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1337_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19182__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09046_ game.CPU.applesa.ab.absxs.body_y\[100\] vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__inv_2
XANTENNA__15586__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold440 game.writer.tracker.frame\[462\] vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09584__B game.CPU.applesa.ab.check_walls.above.walls\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12291__A game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold451 game.writer.tracker.frame\[253\] vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1125_X net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold462 game.writer.tracker.frame\[558\] vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11904__A1 game.CPU.applesa.ab.check_walls.above.walls\[92\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17096__A1 _02491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold473 game.writer.tracker.frame\[278\] vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11904__B2 game.CPU.applesa.ab.check_walls.above.walls\[94\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold484 game.writer.tracker.frame\[50\] vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 game.CPU.applesa.apple_location2_n\[4\] vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11619__B net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout964_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout920 net921 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16843__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout931 _03190_ vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_2
X_09948_ _03196_ _04178_ vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__xnor2_1
Xfanout942 game.CPU.applesa.y\[3\] vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_4
Xfanout953 net957 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__buf_4
XANTENNA_fanout76_A _02690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout964 net973 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__buf_4
XANTENNA__12314__D1 _06101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout975 net976 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_4
Xfanout986 net987 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__buf_2
XANTENNA__17306__B _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout997 net1009 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
X_09879_ _03722_ _03727_ _04032_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__o21a_1
XANTENNA__11194__X _05084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Left_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11910_ net806 net308 _05796_ _05797_ _05285_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_169_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12890_ game.writer.tracker.frame\[62\] game.writer.tracker.frame\[63\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__mux2_1
XANTENNA__14011__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12419__A1_N game.CPU.applesa.ab.absxs.body_x\[35\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09105__A game.CPU.applesa.ab.absxs.body_y\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11841_ game.CPU.applesa.ab.check_walls.above.walls\[150\] net299 _05728_ vssd1 vssd1
+ vccd1 vccd1 _05729_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_200_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14082__A1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14082__B2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17322__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11772_ net571 _05459_ _05659_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__a21oi_1
X_14560_ game.CPU.walls.rand_wall.logic_enable _08426_ _08422_ vssd1 vssd1 vccd1 vccd1
+ _08427_ sky130_fd_sc_hd__a21o_2
XANTENNA__12632__A2 game.CPU.applesa.twoapples.absxs.next_head\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17020__A1 _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13511_ net246 _07382_ _07384_ net190 vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__o31a_1
XANTENNA__14909__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10723_ game.CPU.applesa.ab.absxs.body_y\[39\] _04642_ _04643_ game.CPU.applesa.ab.absxs.body_y\[35\]
+ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__a22o_1
XANTENNA__12466__A game.CPU.applesa.ab.absxs.body_y\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09759__B game.CPU.applesa.ab.check_walls.above.walls\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14909__B2 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14491_ _08206_ _08210_ _08290_ _08364_ _08106_ vssd1 vssd1 vccd1 vccd1 _08365_ sky130_fd_sc_hd__o2111a_1
XANTENNA__11370__A game.CPU.applesa.ab.check_walls.above.walls\[32\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16230_ net162 _02236_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__nand2_8
XFILLER_0_153_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19525__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13442_ net682 _06933_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__or2_1
X_10654_ net1079 _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__nor2_2
XFILLER_0_125_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_190_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_299_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10257__Y _04450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12185__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_298_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11199__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_298_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13373_ net511 _06691_ net702 vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__a21o_1
XFILLER_0_307_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15777__A game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16161_ _02072_ _02074_ _02077_ _02079_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__or4_1
XANTENNA__12753__X _06627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10585_ game.CPU.applesa.ab.absxs.body_x\[112\] _04663_ _04664_ game.CPU.applesa.ab.absxs.body_x\[108\]
+ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__a22o_1
Xclkload18 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload29 clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__inv_6
X_15112_ net1207 net1230 game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1
+ vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__and3_1
X_12324_ net381 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.absxs.next_head\[0\]
+ sky130_fd_sc_hd__inv_2
X_16092_ _03258_ net348 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_310_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13297__A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19920_ clknet_leaf_33_clk game.writer.tracker.next_frame\[515\] net1302 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[515\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19675__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15043_ net1215 net1241 game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1
+ vccd1 vccd1 _00264_ sky130_fd_sc_hd__and3_1
X_12255_ net823 net549 vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17992__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13896__A1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13896__B2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17087__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11206_ _03229_ net319 vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__xnor2_1
X_19851_ clknet_leaf_37_clk game.writer.tracker.next_frame\[446\] net1356 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[446\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_294_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12186_ game.CPU.applesa.ab.check_walls.above.walls\[125\] net547 vssd1 vssd1 vccd1
+ vccd1 _06072_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_71_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11529__B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ game.CPU.applesa.ab.absxs.body_x\[70\] net410 vssd1 vssd1 vccd1 vccd1 _05027_
+ sky130_fd_sc_hd__xnor2_1
X_18802_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[5\] _00539_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[5\] sky130_fd_sc_hd__dfrtp_1
X_19782_ clknet_leaf_24_clk game.writer.tracker.next_frame\[377\] net1344 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[377\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_247_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16401__A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16994_ _02455_ net120 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__and2_1
XFILLER_0_247_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_305_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18733_ clknet_leaf_13_clk _01150_ _00470_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[115\]
+ sky130_fd_sc_hd__dfrtp_4
X_11068_ _03278_ net408 net403 _03349_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__a22o_1
X_15945_ _01953_ _01954_ _01955_ _01956_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_143_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13236__S net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12320__A1 _06142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ net1125 _04226_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__nand2_1
XANTENNA__12320__B2 _06135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15017__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18664_ clknet_leaf_64_clk _01081_ _00401_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[86\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_222_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15876_ game.CPU.applesa.ab.absxs.body_x\[26\] net466 net458 game.CPU.applesa.ab.absxs.body_x\[27\]
+ _01882_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a221o_1
X_17615_ net1973 _03023_ _03025_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__o21a_1
XANTENNA__19055__CLK net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14827_ game.CPU.randy.f1.c1.count\[0\] _04332_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[0\]
+ sky130_fd_sc_hd__and2b_1
XANTENNA__14073__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18595_ clknet_leaf_52_clk _01015_ _00332_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[72\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_203_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14073__B2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18328__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17546_ net1456 _08808_ _02972_ _00293_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14758_ game.CPU.randy.counter1.count1\[17\] _08575_ game.CPU.randy.counter1.count1\[18\]
+ vssd1 vssd1 vccd1 vccd1 _08580_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_290_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13709_ game.writer.tracker.frame\[237\] game.writer.tracker.frame\[239\] game.writer.tracker.frame\[240\]
+ game.writer.tracker.frame\[238\] net968 net998 vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__mux4_1
X_17477_ _02884_ _02899_ _02896_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12376__A game.CPU.applesa.ab.absxs.body_x\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14689_ game.CPU.randy.counter1.count1\[14\] _04347_ _08491_ _08527_ vssd1 vssd1
+ vccd1 vccd1 _08528_ sky130_fd_sc_hd__a31o_1
XFILLER_0_315_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19216_ net1169 _00028_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_possible\[7\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_116_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16428_ _02295_ _02313_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__nand2_2
XFILLER_0_345_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13033__C1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_317_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13584__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19147_ net1188 _00190_ _00818_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[192\]
+ sky130_fd_sc_hd__dfrtp_4
X_16359_ net160 _02342_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__nand2_2
XANTENNA__12663__X _06540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18063__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17314__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10937__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09685__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19078_ net1179 _00114_ _00749_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[123\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16522__B1 _02461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13336__A0 _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11279__X _05169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18029_ net605 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__inv_2
XANTENNA__15876__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17078__A1 _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_285_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout205 net208 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_243_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11362__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout227 net229 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_2
X_09802_ net1155 game.CPU.applesa.ab.check_walls.above.walls\[108\] vssd1 vssd1 vccd1
+ vccd1 _04045_ sky130_fd_sc_hd__xor2_1
XANTENNA__13935__A net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout238 net239 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17407__A _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_238_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout249 net251 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10570__B1 _04594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_340_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09733_ net1136 game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1 _03976_
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout280_A _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16030__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13146__S net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout378_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ net1151 game.CPU.applesa.ab.absxs.body_y\[37\] vssd1 vssd1 vccd1 vccd1 _03907_
+ sky130_fd_sc_hd__or2_1
XANTENNA__17250__A1 _02267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16053__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11174__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09595_ net1092 game.CPU.applesa.ab.absxs.body_x\[74\] vssd1 vssd1 vccd1 vccd1 _03838_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_328_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout166_X net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout545_A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17002__A1 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_254_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11283__D1 _05169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11822__B1 _05689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout712_A _06594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19130__Q game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12286__A game.CPU.applesa.ab.check_walls.above.walls\[135\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09491__A1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1075_X net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17553__A2 _00039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09491__B2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_176_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10518__B _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19698__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1242_X net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09595__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_304_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10370_ net1453 net850 _04195_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_295_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09029_ game.CPU.applesa.ab.absxs.body_x\[27\] vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__inv_2
XANTENNA__10534__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13878__A1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13878__B2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09882__X _04125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12040_ net800 net295 net289 net801 vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a2bb2o_1
Xhold270 game.writer.tracker.frame\[152\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_265_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold281 game.writer.tracker.frame\[84\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 game.writer.tracker.frame\[446\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_X net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_257_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_291_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_187_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16221__A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__B1 _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Left_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout750 net751 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout79_X net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout761 net762 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_129_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout772 game.CPU.applesa.ab.apple_possible\[1\] vssd1 vssd1 vccd1 vccd1 net772
+ sky130_fd_sc_hd__buf_4
XANTENNA__19078__CLK net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout783 game.CPU.applesa.ab.check_walls.above.walls\[183\] vssd1 vssd1 vccd1 vccd1
+ net783 sky130_fd_sc_hd__buf_2
X_13991_ _07858_ _07862_ _07863_ _07864_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_6_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout794 game.CPU.applesa.ab.check_walls.above.walls\[126\] vssd1 vssd1 vccd1 vccd1
+ net794 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11365__A game.CPU.applesa.ab.check_walls.above.walls\[35\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15730_ game.CPU.applesa.ab.absxs.body_x\[15\] net462 vssd1 vssd1 vccd1 vccd1 _01742_
+ sky130_fd_sc_hd__xnor2_1
X_12942_ _06740_ _06743_ net677 vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__mux2_1
XANTENNA__16044__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11084__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15661_ net819 net443 net474 game.CPU.applesa.ab.check_walls.above.walls\[49\] vssd1
+ vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_354_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12895__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ game.writer.tracker.frame\[34\] game.writer.tracker.frame\[35\] net1003 vssd1
+ vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__mux2_1
XANTENNA__13489__S0 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17400_ _04257_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__and2_1
XFILLER_0_358_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14612_ game.CPU.clock1.counter\[9\] _08464_ vssd1 vssd1 vccd1 vccd1 _08465_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_202_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ net600 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__inv_2
X_11824_ game.CPU.applesa.ab.check_walls.above.walls\[127\] net310 vssd1 vssd1 vccd1
+ vccd1 _05712_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15592_ net433 game.CPU.applesa.ab.check_walls.above.walls\[39\] _03397_ net352 vssd1
+ vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_276_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20053__1371 vssd1 vssd1 vccd1 vccd1 _20053__1371/HI net1371 sky130_fd_sc_hd__conb_1
XANTENNA__14395__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17331_ net576 _01449_ _01582_ _08900_ vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__a22o_1
XFILLER_0_200_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10616__A1 game.CPU.applesa.ab.absxs.body_x\[73\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_218_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _03488_ _08414_ vssd1 vssd1 vccd1 vccd1 _08415_ sky130_fd_sc_hd__nor2_1
XANTENNA__17987__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ game.CPU.applesa.ab.check_walls.above.walls\[173\] net306 _05638_ _05641_
+ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__o2111a_1
XANTENNA__18915__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12196__A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Left_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09482__B2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17262_ _02275_ _02309_ _02746_ net1653 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[526\]
+ sky130_fd_sc_hd__a22o_1
X_10706_ game.CPU.applesa.ab.absxs.body_y\[68\] _04625_ _04626_ game.CPU.applesa.ab.absxs.body_y\[64\]
+ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_327_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14474_ _03291_ net1067 net874 game.CPU.applesa.ab.absxs.body_x\[11\] _08346_ vssd1
+ vssd1 vccd1 vccd1 _08348_ sky130_fd_sc_hd__o221a_1
XANTENNA__15003__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11686_ _05571_ _05572_ _05573_ _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__or4_1
XFILLER_0_342_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19001_ net1194 _00228_ _00672_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16213_ _02002_ _02206_ _02218_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__and4_2
X_13425_ _06930_ _06950_ net700 vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__mux2_1
X_17193_ _02501_ net75 _02729_ net1582 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[474\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10637_ net932 game.CPU.applesa.ab.absxs.body_x\[46\] net561 _04686_ vssd1 vssd1
+ vccd1 vccd1 _01117_ sky130_fd_sc_hd__a31o_1
XFILLER_0_314_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13661__S0 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_302_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16144_ game.CPU.applesa.ab.absxs.body_x\[77\] net471 net438 game.CPU.applesa.ab.absxs.body_y\[78\]
+ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__o22a_1
X_13356_ _06659_ _06661_ _06669_ _06660_ net701 net494 vssd1 vssd1 vccd1 vccd1 _07230_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_286_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10568_ _04591_ _04617_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__and2_1
XFILLER_0_178_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_267_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16115__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12307_ game.CPU.applesa.ab.check_walls.above.walls\[189\] net547 vssd1 vssd1 vccd1
+ vccd1 _06193_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_310_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_307_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16075_ _03233_ net471 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__nand2_1
XFILLER_0_310_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13287_ _07115_ _07129_ _07160_ net246 net190 vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__o221a_1
X_10499_ _04358_ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_287_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19903_ clknet_leaf_20_clk game.writer.tracker.next_frame\[498\] net1317 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[498\] sky130_fd_sc_hd__dfrtp_1
X_15026_ net1219 net1248 net819 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__and3_1
XANTENNA__15954__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12238_ _05857_ _06123_ _05855_ _05856_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_229_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10163__B _03527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16807__A1 _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11344__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19834_ clknet_leaf_33_clk game.writer.tracker.next_frame\[429\] net1325 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[429\] sky130_fd_sc_hd__dfrtp_1
X_12169_ game.CPU.applesa.ab.check_walls.above.walls\[158\] net288 net293 net788 vssd1
+ vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_208_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16977_ _02480_ _02634_ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__or2_1
X_19765_ clknet_leaf_29_clk game.writer.tracker.next_frame\[360\] net1291 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[360\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19215__Q game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput5 gpio_in[3] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_265_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15928_ _03446_ net332 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__xnor2_1
X_18716_ clknet_leaf_65_clk _01133_ _00453_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[82\]
+ sky130_fd_sc_hd__dfrtp_4
X_19696_ clknet_leaf_29_clk game.writer.tracker.next_frame\[291\] net1285 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[291\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_274_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18647_ clknet_leaf_12_clk _01064_ _00384_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[53\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_210_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15859_ game.CPU.applesa.ab.absxs.body_x\[115\] net462 vssd1 vssd1 vccd1 vccd1 _01871_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_318_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09380_ net912 game.CPU.applesa.ab.check_walls.above.walls\[8\] _03385_ net1140 _03619_
+ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_160_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18578_ clknet_leaf_61_clk _00998_ _00315_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[35\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15794__A1 game.CPU.applesa.ab.absxs.body_x\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15794__B2 game.CPU.applesa.ab.absxs.body_y\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Left_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17529_ _02782_ net426 _02841_ _02852_ game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1
+ _02957_ sky130_fd_sc_hd__a32o_1
XANTENNA__09399__B game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10619__A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19840__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_318_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16743__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13557__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout126_A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13652__S0 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19990__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12553__B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_329_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13309__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16025__B net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12780__A1 game.writer.tracker.frame\[97\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18521__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1035_A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Left_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11169__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15864__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16312__Y _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19220__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12532__A1 game.CPU.applesa.ab.absxs.body_x\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12532__B2 game.CPU.applesa.ab.absxs.body_y\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09862__B game.CPU.applesa.ab.absxs.body_x\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1202_A game.CPU.walls.rand_wall.good_spot vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout662_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_X clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16976__A _02480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15880__A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09716_ _03952_ _03953_ _03954_ _03958_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_260_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19370__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17223__B2 game.writer.tracker.frame\[497\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18964__Q game.CPU.applesa.ab.check_walls.above.walls\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__A2 game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ net910 game.CPU.applesa.ab.check_walls.above.walls\[152\] game.CPU.applesa.ab.check_walls.above.walls\[153\]
+ net915 vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__o22a_1
XFILLER_0_334_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19878__RESET_B net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14037__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14037__B2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1192_X net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16577__A3 _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13604__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_36_clk_X clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09578_ net923 game.CPU.applesa.ab.check_walls.above.walls\[42\] game.CPU.applesa.ab.check_walls.above.walls\[44\]
+ net895 vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_355_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16982__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_218_Right_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13796__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11632__B net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09837__A2_N game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09464__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11540_ game.CPU.applesa.ab.check_walls.above.walls\[146\] net765 vssd1 vssd1 vccd1
+ vccd1 _05429_ sky130_fd_sc_hd__xor2_2
XFILLER_0_203_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10248__B net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11471_ net827 net261 _05359_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__o21ba_1
XANTENNA__16216__A _06607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_279_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13210_ _07082_ _07083_ net486 vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10422_ game.CPU.up_button.eD1.Q2 game.CPU.up_button.eD1.Q1 vssd1 vssd1 vccd1 vccd1
+ _04567_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_268_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14190_ game.CPU.applesa.ab.absxs.body_y\[99\] net939 vssd1 vssd1 vccd1 vccd1 _08064_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_213_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12463__B net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13141_ game.writer.tracker.frame\[148\] game.writer.tracker.frame\[149\] net1023
+ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__mux2_1
X_10353_ game.CPU.walls.rand_wall.input2 game.CPU.walls.rand_wall.inputa _00290_ vssd1
+ vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__nor3_1
XFILLER_0_150_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13072_ game.writer.tracker.frame\[198\] game.writer.tracker.frame\[199\] net1030
+ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_295_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10284_ net851 game.CPU.applesa.ab.good_spot_next game.CPU.applesa.ab.apple_location\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__a21o_1
XANTENNA__14512__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16900_ net200 _02389_ net92 _02641_ net1911 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[269\]
+ sky130_fd_sc_hd__a32o_1
X_12023_ _05907_ _05908_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__or3_1
XANTENNA__13720__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17880_ net656 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19713__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16831_ net1925 _02610_ _02612_ net132 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[229\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_228_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_302_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19035__Q game.CPU.applesa.ab.check_walls.above.walls\[80\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16598__A1_N net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 net591 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_4
X_19550_ clknet_leaf_34_clk game.writer.tracker.next_frame\[145\] net1328 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[145\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_232_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout591 net625 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_2
XANTENNA__15790__A game.CPU.applesa.ab.absxs.body_x\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16762_ _02419_ net65 net560 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_272_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13974_ net949 game.CPU.applesa.ab.check_walls.above.walls\[86\] vssd1 vssd1 vccd1
+ vccd1 _07848_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_224_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17214__A1 _02533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18501_ net601 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__inv_2
X_15713_ _01721_ _01722_ _01723_ _01724_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__or4_2
X_19481_ clknet_leaf_18_clk game.writer.tracker.next_frame\[76\] net1308 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[76\] sky130_fd_sc_hd__dfrtp_1
X_12925_ net479 _06798_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__or2_1
XFILLER_0_260_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_244_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16693_ _02300_ net61 _02564_ net1579 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[139\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14028__A1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14028__B2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19863__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18432_ net586 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15644_ net813 net445 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_244_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12856_ game.writer.tracker.frame\[300\] game.writer.tracker.frame\[301\] net988
+ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__mux2_1
XANTENNA__19548__RESET_B net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16973__B1 _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_319_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18363_ net597 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__inv_2
X_11807_ net750 _05568_ _05694_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09455__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15575_ game.CPU.kyle.L1.cnt_500hz\[13\] _01587_ game.CPU.kyle.L1.cnt_500hz\[14\]
+ vssd1 vssd1 vccd1 vccd1 game.CPU.en sky130_fd_sc_hd__a21oi_1
XANTENNA__15014__B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12787_ game.writer.tracker.frame\[350\] game.writer.tracker.frame\[351\] net1017
+ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__mux2_1
XANTENNA__09455__B2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17314_ _06701_ net113 _02405_ net733 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__o31a_1
XFILLER_0_260_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14526_ _08369_ _08393_ _08040_ vssd1 vssd1 vccd1 vccd1 _08400_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_185_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11738_ _03463_ net310 vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__xnor2_1
X_18294_ net646 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
XANTENNA__16725__B1 _02577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15949__B net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13539__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_313_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17245_ net175 _02556_ _02742_ game.writer.tracker.frame\[513\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[513\] sky130_fd_sc_hd__a22o_1
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_289_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14457_ game.CPU.applesa.ab.absxs.body_x\[14\] net1056 vssd1 vssd1 vccd1 vccd1 _08331_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11669_ net566 _05551_ _05553_ _05556_ _05557_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_98_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_302_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13408_ net506 _07281_ _07280_ net207 vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__a211o_1
X_17176_ _02311_ _02719_ net557 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11014__B2 net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14388_ _03224_ net1055 net860 game.CPU.applesa.ab.absxs.body_y\[7\] _08260_ vssd1
+ vssd1 vccd1 vccd1 _08262_ sky130_fd_sc_hd__a221o_1
XFILLER_0_330_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16127_ _03249_ net349 net341 _03317_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a22o_1
X_13339_ _07211_ _07212_ net476 vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__mux2_1
XANTENNA__17150__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14503__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16058_ _02061_ _02067_ _02068_ _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__or4b_2
XANTENNA__15684__B net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12514__A1 game.CPU.applesa.ab.absxs.body_x\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16499__C net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15009_ net1221 net1249 net823 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__and3_1
XANTENNA__12514__B2 game.CPU.applesa.ab.absxs.body_y\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16256__A2 _08400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_324_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19817_ clknet_leaf_38_clk game.writer.tracker.next_frame\[412\] net1350 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[412\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_208_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_285_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10621__B _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10113__S _04311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19748_ clknet_leaf_24_clk game.writer.tracker.next_frame\[343\] net1339 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[343\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13475__C1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09501_ net1161 game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1 vccd1
+ vccd1 _03744_ sky130_fd_sc_hd__xor2_1
XANTENNA__10828__A1 net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18784__Q game.CPU.applesa.ab.absxs.body_x\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19971__RESET_B net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14019__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19679_ clknet_leaf_34_clk game.writer.tracker.next_frame\[274\] net1322 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[274\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14019__B2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12829__A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13424__S net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09432_ net907 net796 _03667_ _03671_ _03672_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_338_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16964__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12548__B net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11452__B net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09363_ net920 game.CPU.applesa.ab.check_walls.above.walls\[194\] game.CPU.applesa.ab.check_walls.above.walls\[196\]
+ net891 _03604_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09446__A1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09446__B2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17420__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15519__A1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ net1107 _03423_ net808 net906 vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__o22a_1
XFILLER_0_129_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15859__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_32 _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_43 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09857__B game.CPU.applesa.ab.absxs.body_x\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout410_A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13625__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16036__A game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout508_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout129_X net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_320_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12753__A1 game.writer.tracker.frame\[113\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13947__X _07821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_63_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10764__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18251__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18610__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19736__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12096__A2_N net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15594__B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout877_A net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20052__1370 vssd1 vssd1 vccd1 vccd1 _20052__1370/HI net1370 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_54_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_262_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_273_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09382__B1 game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18760__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19886__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18694__Q game.CPU.applesa.ab.absxs.body_x\[40\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10819__A1 game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_214_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10819__B2 game.CPU.applesa.ab.absxs.body_y\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ net1266 net413 vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12710_ net1057 _06555_ net1048 vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11643__A game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13690_ game.writer.tracker.frame\[511\] net710 net673 game.writer.tracker.frame\[512\]
+ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__o22a_1
XANTENNA__17251__A1_N net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_273_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ _06260_ _06517_ _06261_ _06448_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__or4b_1
XFILLER_0_167_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15360_ _08877_ _08901_ vssd1 vssd1 vccd1 vccd1 _08902_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_16_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12441__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ game.CPU.applesa.ab.absxs.body_x\[16\] net384 vssd1 vssd1 vccd1 vccd1 _06449_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__08952__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14311_ game.CPU.applesa.ab.absxs.body_x\[56\] net1074 vssd1 vssd1 vccd1 vccd1 _08185_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19266__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11523_ game.CPU.applesa.ab.check_walls.above.walls\[40\] net779 vssd1 vssd1 vccd1
+ vccd1 _05412_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_137_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15291_ game.CPU.applesa.twomode.counter_flip game.CPU.applesa.twomode.number\[4\]
+ vssd1 vssd1 vccd1 vccd1 _08841_ sky130_fd_sc_hd__and2b_1
XANTENNA__13616__S0 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17030_ _02370_ _02670_ net717 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14242_ _08111_ _08112_ _08113_ vssd1 vssd1 vccd1 vccd1 _08116_ sky130_fd_sc_hd__or3_1
XFILLER_0_150_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11454_ net812 net257 net316 net813 vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12193__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ _04341_ _04349_ game.CPU.randy.f1.state\[2\] vssd1 vssd1 vccd1 vccd1 _04553_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__15785__A game.CPU.applesa.ab.absxs.body_y\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14173_ game.CPU.applesa.ab.absxs.body_y\[106\] net953 vssd1 vssd1 vccd1 vccd1 _08047_
+ sky130_fd_sc_hd__xor2_1
X_11385_ net784 net251 _05273_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__a21oi_1
X_13124_ _06994_ _06996_ net696 vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__mux2_1
X_10336_ game.CPU.randy.f1.a1.count\[5\] _04489_ game.CPU.randy.f1.a1.count\[6\] vssd1
+ vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__a21o_1
X_18981_ net1197 _00206_ _00652_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_284_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13055_ net492 _06928_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__or2_1
X_17932_ net660 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__inv_2
X_10267_ net766 net742 vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_226_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1320 net1323 vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16238__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ net786 net294 net289 game.CPU.applesa.ab.check_walls.above.walls\[166\] vssd1
+ vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__a22o_1
XANTENNA__09373__B1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1331 net1332 vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__buf_2
X_17863_ net833 _03173_ _03147_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__o21ai_1
Xfanout1342 net1343 vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__clkbuf_4
X_10198_ net1168 net759 vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__nand2_1
XANTENNA__15009__B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1353 net1359 vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__buf_2
XANTENNA__16789__A3 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15446__B1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19602_ clknet_leaf_22_clk game.writer.tracker.next_frame\[197\] net1342 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[197\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16814_ _02503_ net105 _02604_ net1865 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[220\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13457__C1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17794_ net883 _03134_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19533_ clknet_leaf_23_clk game.writer.tracker.next_frame\[128\] net1344 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[128\] sky130_fd_sc_hd__dfrtp_1
X_16745_ game.writer.tracker.frame\[172\] _02583_ vssd1 vssd1 vccd1 vccd1 _02584_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_198_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13957_ _07827_ _07828_ _07829_ _07830_ vssd1 vssd1 vccd1 vccd1 _07831_ sky130_fd_sc_hd__or4_1
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19464_ clknet_leaf_40_clk game.writer.tracker.next_frame\[59\] net1354 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[59\] sky130_fd_sc_hd__dfrtp_1
X_12908_ game.writer.tracker.frame\[54\] game.writer.tracker.frame\[55\] net1037 vssd1
+ vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__mux2_1
XANTENNA__11483__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15025__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16676_ game.writer.tracker.frame\[129\] _02554_ _02557_ vssd1 vssd1 vccd1 vccd1
+ game.writer.tracker.next_frame\[129\] sky130_fd_sc_hd__a21o_1
XFILLER_0_186_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_319_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13888_ net950 game.CPU.applesa.ab.check_walls.above.walls\[102\] vssd1 vssd1 vccd1
+ vccd1 _07762_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12368__B net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_295_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15627_ _03480_ net350 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__xnor2_1
X_18415_ net626 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__inv_2
X_12839_ _06711_ _06712_ net510 vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__mux2_1
XANTENNA__19609__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19395_ clknet_leaf_55_clk net2 net1280 vssd1 vssd1 vccd1 vccd1 game.writer.control.button5.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09428__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_237_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09428__B2 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16408__X _02378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18336__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10038__A2 _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18346_ net594 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__inv_2
XANTENNA__09958__A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15558_ _01571_ _01577_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__nand2_2
XFILLER_0_185_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16159__D1 _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15679__B net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12983__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14509_ game.CPU.apple_location2\[6\] net947 vssd1 vssd1 vccd1 vccd1 _08383_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18277_ net641 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
XANTENNA__09677__B game.CPU.applesa.ab.absxs.body_x\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15489_ _08368_ _08394_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13607__S0 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17228_ _02413_ _02720_ net727 vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__o21a_1
XANTENNA__18633__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14185__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19759__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17159_ _02237_ net122 vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__nand2_2
XFILLER_0_12_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09600__B2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_326_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09693__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09981_ game.CPU.applesa.off_bc.Q2 game.CPU.applesa.off_bc.Q1 vssd1 vssd1 vccd1 vccd1
+ _04207_ sky130_fd_sc_hd__and2b_4
XANTENNA__13927__B game.CPU.applesa.ab.check_walls.above.walls\[34\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16303__B _02301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload28_A clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18783__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14104__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11447__B net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17415__A _02779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19139__CLK net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout360_A net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_315_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout458_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11463__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_337_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12278__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11182__B net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09415_ net1136 game.CPU.applesa.ab.absxs.body_y\[98\] vssd1 vssd1 vccd1 vccd1 _03658_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_149_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout246_X net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A _08799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18246__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14412__B2 game.CPU.applesa.ab.absxs.body_y\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_325_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09868__A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12423__B1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ net1142 game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1 _03589_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_353_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17301__C_N _02379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09277_ net758 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_306_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1155_X net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14176__B1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout994_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_348_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12821__S1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11170_ net1267 net324 vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_132_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_274_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14479__B2 game.CPU.applesa.ab.absxs.body_y\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10121_ _04320_ game.CPU.applesa.apple_location2_n\[0\] _04311_ vssd1 vssd1 vccd1
+ vccd1 _01340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11638__A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14014__A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13151__A1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__A game.CPU.applesa.ab.absxs.body_y\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ game.CPU.applesa.twoapples.count_luck\[7\] game.CPU.applesa.twoapples.count_luck\[5\]
+ game.CPU.applesa.twoapples.count_luck\[6\] vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__or3b_1
XFILLER_0_274_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11357__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ net1561 _08649_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[13\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_242_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13811_ game.writer.tracker.frame\[413\] game.writer.tracker.frame\[415\] game.writer.tracker.frame\[416\]
+ game.writer.tracker.frame\[414\] net980 net1037 vssd1 vssd1 vccd1 vccd1 _07685_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_230_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14791_ game.CPU.randy.counter1.count\[5\] game.CPU.randy.counter1.count\[4\] _08604_
+ vssd1 vssd1 vccd1 vccd1 _08608_ sky130_fd_sc_hd__and3_1
XANTENNA__09658__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_221_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09658__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_270_Right_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_230_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16530_ _02298_ _02340_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__nor2_8
XFILLER_0_225_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_329_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13742_ _07614_ _07615_ net491 vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__mux2_1
XANTENNA__16928__B1 _02650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12662__B1 _06538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ _04837_ _04838_ _04842_ _04843_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__or4_1
XANTENNA__16883__B _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17196__A3 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__B net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16461_ net169 net112 net69 _02414_ net1778 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[55\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13673_ game.writer.tracker.frame\[457\] game.writer.tracker.frame\[459\] game.writer.tracker.frame\[460\]
+ game.writer.tracker.frame\[458\] net974 net1013 vssd1 vssd1 vccd1 vccd1 _07547_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_317_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10885_ net1171 net547 net551 game.CPU.applesa.ab.YMAX\[0\] vssd1 vssd1 vccd1 vccd1
+ _04787_ sky130_fd_sc_hd__o211a_1
XFILLER_0_356_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13837__S0 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18200_ net580 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__inv_2
XANTENNA__15600__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15412_ _03366_ _08939_ _01439_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_344_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18656__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09778__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12624_ _06364_ _06365_ _06366_ _06367_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__or4_1
X_19180_ clknet_leaf_6_clk _01299_ _00842_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_16392_ net1941 net721 _02366_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[36\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__19901__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11768__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18131_ net578 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15343_ game.writer.updater.commands.cmd_num\[1\] _08878_ _08880_ _08884_ vssd1 vssd1
+ vccd1 vccd1 _08885_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12555_ game.CPU.applesa.ab.absxs.body_x\[84\] net381 vssd1 vssd1 vccd1 vccd1 _06432_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09497__B game.CPU.applesa.ab.check_walls.above.walls\[48\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09830__A1 net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09830__B2 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_310_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18062_ net613 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__inv_2
X_11506_ net831 net262 vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__nand2_1
X_15274_ _08817_ _01261_ vssd1 vssd1 vccd1 vccd1 _08828_ sky130_fd_sc_hd__nand2_1
XFILLER_0_324_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12486_ game.CPU.applesa.ab.absxs.body_y\[82\] net517 vssd1 vssd1 vccd1 vccd1 _06363_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__15011__C game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19983__Q game.CPU.applesa.y\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17013_ _02503_ net89 _02675_ net1606 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[348\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_232_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14225_ game.CPU.applesa.ab.absxs.body_x\[42\] net1059 vssd1 vssd1 vccd1 vccd1 _08099_
+ sky130_fd_sc_hd__or2_1
X_11437_ net746 _05321_ _05325_ _05315_ _05316_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_111_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16404__A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14156_ net904 net853 vssd1 vssd1 vccd1 vccd1 _08030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11368_ game.CPU.applesa.ab.check_walls.above.walls\[33\] net771 vssd1 vssd1 vccd1
+ vccd1 _05257_ sky130_fd_sc_hd__xor2_1
XFILLER_0_265_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ net511 _06927_ _06929_ net228 vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__o211a_1
XANTENNA__10743__A3 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ game.CPU.randy.f1.a1.count\[10\] net740 _04493_ vssd1 vssd1 vccd1 vccd1 _04500_
+ sky130_fd_sc_hd__and3_1
X_18964_ net1199 _00287_ _00635_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_14087_ net1073 _03427_ _03430_ net952 _07960_ vssd1 vssd1 vccd1 vccd1 _07961_ sky130_fd_sc_hd__a221o_1
X_11299_ _04876_ _04878_ _05188_ _05127_ _05044_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__o311a_1
XFILLER_0_237_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12556__A2_N net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13038_ _06869_ _06884_ net699 vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__mux2_1
X_17915_ net607 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__inv_2
XANTENNA__09018__A game.CPU.applesa.ab.absxs.body_x\[73\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09897__A1 _03812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18895_ clknet_leaf_1_clk _00000_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_146_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13693__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16410__Y _02379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1150 net1151 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_321_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1161 game.CPU.applesa.ab.snake_head_y\[0\] vssd1 vssd1 vccd1 vccd1 net1161
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__19563__RESET_B net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17846_ _03155_ _03170_ _03171_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__and3_1
XFILLER_0_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1172 net1173 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__clkbuf_4
Xfanout1183 net1184 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__buf_2
Xfanout1194 net1195 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_206_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19431__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14989_ net1227 net1254 game.CPU.applesa.ab.check_walls.above.walls\[17\] vssd1 vssd1
+ vccd1 vccd1 _00205_ sky130_fd_sc_hd__and3_1
X_17777_ game.CPU.applesa.twoapples.count\[2\] game.CPU.applesa.twoapples.count\[1\]
+ _03125_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__nand3_1
XFILLER_0_345_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19516_ clknet_leaf_28_clk game.writer.tracker.next_frame\[111\] net1287 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[111\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10259__A2 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16728_ net160 net56 net106 _02578_ net1807 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[160\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_18_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12653__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16919__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13850__C1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16659_ net153 net128 _02423_ _02546_ net1549 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[122\]
+ sky130_fd_sc_hd__a32o_1
X_19447_ clknet_leaf_47_clk game.writer.tracker.next_frame\[42\] net1298 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[42\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20043__1367 vssd1 vssd1 vccd1 vccd1 _20043__1367/HI net1367 sky130_fd_sc_hd__conb_1
XANTENNA__16138__X _02150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09200_ net793 vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__inv_2
XANTENNA__09688__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19581__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19378_ clknet_leaf_4_clk _01384_ _00959_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.snake_head_y\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_335_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11759__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_323_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10416__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09131_ game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1 vccd1
+ _03380_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_332_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18329_ net599 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__inv_2
XANTENNA__11730__B net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09062_ game.CPU.applesa.ab.absxs.body_y\[44\] vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16698__A2 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_301_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold600 game.CPU.clock1.counter\[19\] vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout206_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold611 game.CPU.applesa.ab.apple_location\[3\] vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10719__B1 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold622 game.writer.tracker.frame\[128\] vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13381__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold633 game.writer.tracker.frame\[549\] vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 game.writer.tracker.frame\[554\] vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold655 game.writer.tracker.frame\[125\] vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17111__A3 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold666 game.writer.updater.commands.count\[4\] vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16033__B net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11458__A game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10362__A game.CPU.walls.rand_wall.input2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ net1128 _04193_ net754 vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_176_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11177__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14330__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16870__A2 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15872__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _03830_ _03835_ _03903_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout196_X net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_181_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12892__A0 _06762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout742_A _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_358_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19133__Q game.CPU.applesa.ab.check_walls.above.walls\[178\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12289__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18679__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19924__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_257_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_342_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout530_X net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13819__S0 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13612__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_270_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_342_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10670_ _04595_ _04655_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__nor2_2
XFILLER_0_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12947__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09329_ net925 game.CPU.applesa.ab.absxs.body_x\[83\] game.CPU.applesa.ab.absxs.body_y\[83\]
+ net906 vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_63_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14149__B1 _07821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12340_ _04257_ _06217_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout997_X net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12271_ _06154_ _06155_ _06156_ _06153_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__or4b_1
XFILLER_0_287_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14010_ _07877_ _07878_ _07879_ _07883_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__or4_1
XANTENNA__12175__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11222_ _03313_ net534 vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_268_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15649__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__A game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11153_ _05033_ _05037_ _05042_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_281_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16310__B2 _08028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13124__A1 _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ _04252_ _04258_ _04310_ _04256_ _03492_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__o221ai_4
XANTENNA__16861__A2 _02413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15961_ _03391_ net351 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11087__B net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084_ game.CPU.applesa.ab.absxs.body_y\[61\] net542 vssd1 vssd1 vccd1 vccd1 _04974_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__15782__B net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12898__S net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18796__D _00039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_297_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16230__Y _02238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19454__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13675__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14912_ game.CPU.applesa.ab.XMAX\[0\] _08414_ _08417_ game.CPU.applesa.ab.XMAX\[1\]
+ vssd1 vssd1 vccd1 vccd1 _08689_ sky130_fd_sc_hd__a22o_1
X_10035_ game.CPU.applesa.ab.XMAX\[1\] _04210_ _04212_ game.CPU.applesa.ab.XMAX\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__a22o_1
X_17700_ game.CPU.walls.rand_wall.count\[2\] game.CPU.walls.rand_wall.count\[1\] _03075_
+ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__nand3_1
XANTENNA__09780__B net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18680_ clknet_leaf_13_clk _01097_ _00417_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[118\]
+ sky130_fd_sc_hd__dfrtp_4
X_15892_ game.CPU.applesa.ab.absxs.body_x\[40\] net273 vssd1 vssd1 vccd1 vccd1 _01904_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__14398__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17631_ _03035_ net429 _03034_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__and3b_1
X_14843_ game.CPU.randy.f1.c1.count\[6\] _08638_ vssd1 vssd1 vccd1 vccd1 _08641_ sky130_fd_sc_hd__nand2_1
XFILLER_0_349_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_357_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15821__B1 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17562_ net740 _02851_ _02952_ _02848_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__a22o_1
XANTENNA__11438__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14774_ game.CPU.randy.counter1.count\[15\] net265 _08582_ _08594_ vssd1 vssd1 vccd1
+ vccd1 _08595_ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11438__B2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11986_ _05265_ _05270_ _05872_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__or3_1
XANTENNA__15006__C game.CPU.applesa.ab.check_walls.above.walls\[34\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16513_ _02240_ net159 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__nor2_4
X_19301_ clknet_leaf_56_clk game.CPU.applesa.ab.check_walls.below.collision _00916_
+ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.collision_down sky130_fd_sc_hd__dfrtp_1
X_13725_ net511 _07594_ _07595_ _07598_ net228 vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__a311o_2
XTAP_TAPCELL_ROW_15_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16377__A1 game.writer.tracker.frame\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_230_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ game.CPU.applesa.ab.absxs.body_x\[10\] net409 net398 game.CPU.applesa.ab.absxs.body_y\[11\]
+ _04818_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__a221o_1
X_17493_ game.CPU.speed1.Qa\[1\] _02782_ net427 _02921_ vssd1 vssd1 vccd1 vccd1 _02922_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_357_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_292_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16371__C_N _02351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16444_ net1869 _02395_ _02404_ net112 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[50\]
+ sky130_fd_sc_hd__a22o_1
X_19232_ clknet_leaf_57_clk net1423 _00870_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.normal1.number\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__14388__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13656_ _07528_ _07529_ net481 vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__mux2_1
XANTENNA__10661__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_234_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10868_ _04741_ _04742_ _04756_ _04770_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__or4_1
XFILLER_0_344_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12938__A1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16118__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_305_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12607_ _06377_ _06378_ _06381_ _06483_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__or4b_1
X_19163_ clknet_leaf_67_clk _01283_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count_luck\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16375_ net198 _02353_ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__nor2_2
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15022__B net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13587_ _07459_ _07460_ net510 vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10949__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10799_ game.CPU.applesa.ab.absxs.body_y\[34\] _04696_ _04697_ game.CPU.applesa.ab.absxs.body_y\[30\]
+ vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__a22o_1
X_18114_ net584 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15326_ game.CPU.applesa.twomode.number\[6\] _08864_ vssd1 vssd1 vccd1 vccd1 _08870_
+ sky130_fd_sc_hd__nor2_1
X_19094_ net1177 _00131_ _00765_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[139\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12480__A2_N net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12538_ game.CPU.applesa.ab.absxs.body_x\[40\] net384 _06413_ _06414_ vssd1 vssd1
+ vccd1 vccd1 _06415_ sky130_fd_sc_hd__a211o_1
XANTENNA__15957__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18045_ net659 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__inv_2
XFILLER_0_312_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15257_ _08812_ _08814_ vssd1 vssd1 vccd1 vccd1 _08815_ sky130_fd_sc_hd__nor2_1
X_12469_ game.CPU.applesa.ab.absxs.body_x\[13\] net378 net366 game.CPU.applesa.ab.absxs.body_y\[15\]
+ _06342_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__o221a_1
XFILLER_0_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_340_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13110__X _06984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09567__B1 game.CPU.applesa.ab.absxs.body_y\[76\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14208_ _03230_ net1061 net855 game.CPU.applesa.ab.absxs.body_y\[94\] vssd1 vssd1
+ vccd1 vccd1 _08082_ sky130_fd_sc_hd__a22o_1
XANTENNA__13869__A2_N net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10177__A1 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15188_ _08761_ _08762_ vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14139_ _08009_ _08010_ _08011_ _08012_ vssd1 vssd1 vccd1 vccd1 _08013_ sky130_fd_sc_hd__or4_1
XANTENNA__16301__A1 _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout409 net410 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16421__X _02387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19996_ clknet_leaf_45_clk _01420_ net1304 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11709__C _05566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14312__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16852__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18947_ clknet_leaf_68_clk _00076_ _00618_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15692__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09680_ net1111 game.CPU.applesa.ab.absxs.body_x\[100\] vssd1 vssd1 vccd1 vccd1 _03923_
+ sky130_fd_sc_hd__or2_1
XANTENNA__10910__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18878_ clknet_leaf_5_clk game.CPU.randy.f1.c1.innerCount\[8\] _00573_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16300__C _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19947__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17829_ game.writer.updater.commands.count\[3\] _03153_ game.writer.updater.commands.count\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__a21o_1
XANTENNA__10885__C1 game.CPU.applesa.ab.YMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14076__C1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15812__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10121__S _04311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13823__C1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_334_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13940__B game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16309__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout156_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_308_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11460__B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1065_A net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09114_ game.writer.updater.commands.mode\[2\] vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__inv_2
XANTENNA__19327__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13029__S1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09045_ game.CPU.applesa.ab.absxs.body_y\[101\] vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout111_X net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1232_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12572__A game.CPU.applesa.ab.absxs.body_x\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_288_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14490__C _08363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_345_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold430 game.writer.tracker.frame\[397\] vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold441 game.writer.tracker.frame\[318\] vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12291__B net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 game.writer.tracker.frame\[61\] vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A _06600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19128__Q game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold463 game.writer.tracker.frame\[349\] vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19477__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11904__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17096__A2 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold474 game.writer.tracker.frame\[118\] vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 game.writer.tracker.frame\[351\] vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13106__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold496 game.writer.tracker.frame\[281\] vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout910 net913 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_8
Xfanout921 _03193_ vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_8
XANTENNA__14303__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16843__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18967__Q game.CPU.applesa.ab.check_walls.above.walls\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout932 net937 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_4
X_09947_ _04179_ _04182_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout943 net944 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__buf_4
Xfanout954 net955 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout957_A game.CPU.applesa.y\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net973 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_4
Xfanout976 net977 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11668__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ _03806_ _03950_ _03992_ _04075_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__and4_2
Xfanout987 net1042 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__clkbuf_8
XANTENNA__17306__C _02394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout998 net1000 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16056__B1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout69_A _02331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11012__A2_N net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_224_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11840_ _05427_ _05725_ _05726_ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__or4_1
XFILLER_0_197_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19798__Q game.writer.tracker.frame\[393\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_339_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17322__B _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11771_ net747 _05460_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout912_X net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16219__A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13510_ net202 _07300_ _07383_ net277 vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__o211a_1
XANTENNA__11651__A game.CPU.applesa.ab.check_walls.above.walls\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17020__A2 _02670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10722_ game.CPU.applesa.ab.absxs.body_y\[44\] _04640_ _04641_ game.CPU.applesa.ab.absxs.body_y\[40\]
+ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__a22o_1
X_14490_ _08092_ _08311_ _08363_ vssd1 vssd1 vccd1 vccd1 _08364_ sky130_fd_sc_hd__and3_1
XFILLER_0_165_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12573__A1_N game.CPU.applesa.ab.absxs.body_y\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12466__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09121__A game.CPU.applesa.ab.XMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13441_ _07313_ _07314_ net492 vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__mux2_1
XANTENNA__11370__B net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10653_ _04174_ _04695_ _04642_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_190_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16160_ _02164_ _02167_ _02168_ _02169_ _02171_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__o221a_1
XFILLER_0_106_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13372_ _07242_ _07245_ net220 vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__mux2_1
XANTENNA__15777__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ game.CPU.applesa.ab.absxs.body_x\[113\] _04663_ _04664_ game.CPU.applesa.ab.absxs.body_x\[109\]
+ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_101_Left_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16225__Y _02233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload19 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__inv_16
X_15111_ net1204 net1230 game.CPU.applesa.ab.check_walls.above.walls\[139\] vssd1
+ vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12323_ _04212_ _04258_ _04808_ net1162 vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16091_ game.CPU.applesa.ab.absxs.body_y\[110\] net441 vssd1 vssd1 vccd1 vccd1 _02103_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__16531__A1 net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_322_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09549__B1 game.CPU.applesa.ab.absxs.body_y\[113\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12779__S0 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15042_ net1219 net1248 net814 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__and3_1
XFILLER_0_294_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12254_ net802 net423 vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19038__Q game.CPU.applesa.ab.check_walls.above.walls\[83\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13896__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ game.CPU.applesa.ab.absxs.body_x\[92\] net326 vssd1 vssd1 vccd1 vccd1 _05095_
+ sky130_fd_sc_hd__or2_1
XANTENNA__15793__A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19850_ clknet_leaf_40_clk game.writer.tracker.next_frame\[445\] net1356 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[445\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17087__A2 _02393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12185_ net816 net423 vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_208_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20042__1366 vssd1 vssd1 vccd1 vccd1 _20042__1366/HI net1366 sky130_fd_sc_hd__conb_1
X_18801_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[4\] _00538_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[4\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09791__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ game.CPU.applesa.ab.absxs.body_x\[68\] net325 vssd1 vssd1 vccd1 vccd1 _05026_
+ sky130_fd_sc_hd__or2_1
X_19781_ clknet_leaf_23_clk game.writer.tracker.next_frame\[376\] net1344 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[376\] sky130_fd_sc_hd__dfrtp_2
X_16993_ _02476_ net88 _02668_ net1773 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[335\]
+ sky130_fd_sc_hd__a22o_1
X_18732_ clknet_leaf_13_clk _01149_ _00469_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[114\]
+ sky130_fd_sc_hd__dfrtp_4
X_11067_ game.CPU.applesa.ab.absxs.body_x\[26\] net411 vssd1 vssd1 vccd1 vccd1 _04957_
+ sky130_fd_sc_hd__nor2_1
X_15944_ _03405_ game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 _01956_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_143_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ net1163 game.CPU.applesa.out_random_2\[7\] vssd1 vssd1 vccd1 vccd1 _04226_
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_188_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18663_ clknet_leaf_64_clk _01080_ _00400_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[85\]
+ sky130_fd_sc_hd__dfrtp_4
X_15875_ _03279_ net347 net340 _03350_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a22o_1
XANTENNA__15017__B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16598__B2 _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_240_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ net139 _08630_ vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__and2_1
X_17614_ game.CPU.kyle.L1.cnt_20ms\[10\] _03023_ net577 vssd1 vssd1 vccd1 vccd1 _03025_
+ sky130_fd_sc_hd__a21oi_1
X_18594_ clknet_leaf_50_clk _01014_ _00331_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[67\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14073__A2 game.CPU.applesa.ab.check_walls.above.walls\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17545_ _04612_ _02939_ _02963_ _02971_ _02879_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__a2111o_1
X_14757_ _03495_ _03496_ _08575_ vssd1 vssd1 vccd1 vccd1 _08579_ sky130_fd_sc_hd__or3b_1
X_11969_ game.CPU.applesa.ab.check_walls.above.walls\[148\] net551 vssd1 vssd1 vccd1
+ vccd1 _05856_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_82_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13252__S net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17011__A2 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ net241 _07573_ _07581_ net177 _07563_ vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__o311a_1
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11831__A1 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17476_ _02901_ _02902_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__nand2_1
XANTENNA__11292__C1 _05105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14688_ game.CPU.randy.counter1.count1\[15\] _08499_ _08526_ vssd1 vssd1 vccd1 vccd1
+ _08527_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_317_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12376__B net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19215_ net1169 _00027_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_possible\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_132_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13639_ _07508_ _07512_ net215 vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__mux2_1
X_16427_ net115 _02310_ net164 _02388_ net1681 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[46\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_73_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_345_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11797__A1_N net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16358_ net197 _02301_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__nor2_2
X_19146_ net1187 _00189_ _00817_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[191\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15687__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17314__A3 _02405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15309_ game.CPU.applesa.twomode.number\[7\] _08851_ vssd1 vssd1 vccd1 vccd1 _08856_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16289_ net222 net235 net195 _02290_ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__or4_4
X_19077_ net1179 _00113_ _00748_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[122\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09685__B net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16522__B2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18028_ net662 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17078__A2 _02693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16151__X _02163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11898__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11898__B2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout206 net208 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_8
Xfanout217 net218 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
X_09801_ net907 net800 game.CPU.applesa.ab.check_walls.above.walls\[106\] net921 vssd1
+ vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__a2bb2o_1
Xfanout228 net229 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_4
XFILLER_0_226_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13935__B net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19979_ clknet_leaf_42_clk game.writer.tracker.next_frame\[574\] net1326 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[574\] sky130_fd_sc_hd__dfrtp_1
Xfanout239 net243 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkload10_A clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10570__A1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13427__S net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15990__X _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11295__X _05185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ net1136 game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1 _03975_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_340_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09206__A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09663_ net1148 game.CPU.applesa.ab.absxs.body_y\[37\] vssd1 vssd1 vccd1 vccd1 _03906_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__16589__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout273_A game.CPU.walls.rand_wall.abduyd.next_wall\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17250__A2 _02275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09594_ net1092 game.CPU.applesa.ab.absxs.body_x\[74\] vssd1 vssd1 vccd1 vccd1 _03837_
+ sky130_fd_sc_hd__or2_1
XANTENNA__13272__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout440_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16039__A game.CPU.applesa.ab.absxs.body_x\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1182_A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout159_X net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_254_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10625__A2 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16210__B1 _02221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_336_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16761__A1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18254__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1068_X net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12378__A2 game.CPU.applesa.twoapples.absxs.next_head\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15597__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10389__B2 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17305__A3 _02390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10928__A3 game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09595__B game.CPU.applesa.ab.absxs.body_x\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1235_X net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09028_ game.CPU.applesa.ab.absxs.body_x\[32\] vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10534__B _04639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold260 game.writer.tracker.frame\[383\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold271 game.writer.tracker.frame\[369\] vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_265_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold282 game.writer.tracker.frame\[529\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_348_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold293 game.writer.tracker.frame\[286\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_207_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16816__A2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_257_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_284_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_187_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10561__A1 game.CPU.applesa.ab.absxs.body_x\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16221__B net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 net741 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_2
XANTENNA__10561__B2 game.CPU.applesa.ab.absxs.body_x\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13337__S net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout751 _04442_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_4
XANTENNA__11646__A game.CPU.applesa.ab.check_walls.above.walls\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout762 net764 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_129_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14022__A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout773 net774 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__buf_4
X_13990_ net890 game.CPU.applesa.ab.check_walls.above.walls\[16\] game.CPU.applesa.ab.check_walls.above.walls\[18\]
+ net879 _07860_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_6_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16029__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout784 game.CPU.applesa.ab.check_walls.above.walls\[180\] vssd1 vssd1 vccd1 vccd1
+ net784 sky130_fd_sc_hd__buf_2
Xfanout795 game.CPU.applesa.ab.check_walls.above.walls\[125\] vssd1 vssd1 vccd1 vccd1
+ net795 sky130_fd_sc_hd__clkbuf_4
X_12941_ net500 _06814_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11365__B net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17241__A2 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15660_ _03407_ net349 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__xnor2_1
X_12872_ game.writer.tracker.frame\[38\] game.writer.tracker.frame\[39\] net1003 vssd1
+ vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_354_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _08464_ net268 _08463_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[8\]
+ sky130_fd_sc_hd__and3b_1
X_11823_ _05655_ _05663_ _05671_ _05710_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__or4b_1
XANTENNA__13263__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ game.CPU.applesa.ab.check_walls.above.walls\[34\] net467 vssd1 vssd1 vccd1
+ vccd1 _01603_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12477__A game.CPU.applesa.ab.absxs.body_x\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13802__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_276_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17330_ _08916_ _01454_ _08937_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__mux2_1
XANTENNA__11381__A game.CPU.applesa.ab.check_walls.above.walls\[176\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14542_ net1176 game.CPU.walls.abc.number_out\[0\] vssd1 vssd1 vccd1 vccd1 _08414_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_339_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10616__A2 _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11754_ net785 net391 net306 game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1
+ vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11813__A1 game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_218_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12196__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17261_ net207 net112 _02389_ _02746_ net1879 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[525\]
+ sky130_fd_sc_hd__a32o_1
X_10705_ game.CPU.applesa.ab.absxs.body_y\[69\] _04625_ _04626_ game.CPU.applesa.ab.absxs.body_y\[65\]
+ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__a22o_1
XANTENNA__15788__A game.CPU.applesa.ab.absxs.body_x\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14473_ _03292_ net1074 net858 game.CPU.applesa.ab.absxs.body_y\[11\] vssd1 vssd1
+ vccd1 vccd1 _08347_ sky130_fd_sc_hd__a22o_1
XANTENNA__19642__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11685_ net567 _05569_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_299_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16752__B2 game.writer.tracker.frame\[176\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_327_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16212_ _01931_ _01934_ _01939_ _02223_ _01814_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__o311a_2
XFILLER_0_102_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19000_ net1194 _00227_ _00671_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[45\]
+ sky130_fd_sc_hd__dfrtp_4
X_13424_ _06949_ _06951_ net693 vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09786__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_342_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17192_ _02499_ net74 net558 vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a21oi_1
X_10636_ _03272_ net561 vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15820__A2_N net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13661__S1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16143_ net1267 net356 net335 _03300_ _01860_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__o221a_1
XFILLER_0_342_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13355_ _07224_ _07225_ _07228_ net278 net246 vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10567_ game.CPU.applesa.ab.absxs.body_x\[12\] _04653_ _04654_ game.CPU.applesa.ab.absxs.body_x\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__a22o_1
XANTENNA__13318__A1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14515__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ _06188_ _06189_ _06190_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__or4_1
XANTENNA__19792__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16074_ game.CPU.applesa.ab.absxs.body_x\[85\] net350 vssd1 vssd1 vccd1 vccd1 _02086_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_307_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13286_ _07142_ _07143_ _07151_ _07159_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__o22a_1
XFILLER_0_267_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10498_ net1122 _04579_ _04584_ _04619_ _04620_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__o311a_1
XANTENNA__13595__X _07469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_287_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19902_ clknet_leaf_28_clk game.writer.tracker.next_frame\[497\] net1288 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[497\] sky130_fd_sc_hd__dfrtp_1
X_15025_ net1221 net1249 game.CPU.applesa.ab.check_walls.above.walls\[53\] vssd1 vssd1
+ vccd1 vccd1 _00245_ sky130_fd_sc_hd__and3_1
XFILLER_0_258_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12237_ game.CPU.applesa.ab.check_walls.above.walls\[149\] net547 vssd1 vssd1 vccd1
+ vccd1 _06123_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16412__A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_229_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12541__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16807__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19833_ clknet_leaf_33_clk game.writer.tracker.next_frame\[428\] net1325 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[428\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_258_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_248_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12168_ _06052_ _06053_ _06054_ _06051_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__a211o_1
XANTENNA__19022__CLK net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10552__B2 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11119_ game.CPU.applesa.ab.absxs.body_x\[19\] net407 vssd1 vssd1 vccd1 vccd1 _05009_
+ sky130_fd_sc_hd__nand2_1
X_19764_ clknet_leaf_30_clk game.writer.tracker.next_frame\[359\] net1292 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[359\] sky130_fd_sc_hd__dfrtp_1
X_16976_ _02480_ _02634_ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__nor2_1
XFILLER_0_223_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11549__A2_N net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12099_ net798 net387 vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__nand2_1
XFILLER_0_290_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14294__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18715_ clknet_leaf_65_clk _01132_ _00452_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[81\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09026__A game.CPU.applesa.ab.absxs.body_x\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15970__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15927_ _01923_ _01924_ _01927_ _01928_ _01938_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__a221o_1
Xinput6 gpio_in[4] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12939__X _06813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19695_ clknet_leaf_29_clk game.writer.tracker.next_frame\[290\] net1285 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[290\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11843__X _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_349_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17232__A2 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18646_ clknet_leaf_12_clk _01063_ _00383_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[52\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__19172__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15858_ _01865_ _01867_ _01868_ _01869_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__or4_1
XFILLER_0_349_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_318_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14809_ game.CPU.randy.counter1.count\[10\] game.CPU.randy.counter1.count\[9\] _08614_
+ game.CPU.randy.counter1.count\[11\] vssd1 vssd1 vccd1 vccd1 _08620_ sky130_fd_sc_hd__a31o_1
XFILLER_0_176_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18577_ clknet_leaf_58_clk _00997_ _00314_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[34\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12387__A game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10459__X _04594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15789_ game.CPU.applesa.ab.absxs.body_y\[72\] net454 vssd1 vssd1 vccd1 vccd1 _01801_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__15794__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17528_ _03218_ _04257_ net428 _02954_ _02955_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__a311o_1
XFILLER_0_290_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16743__A1 _02379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17459_ net1116 _04638_ _02784_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18074__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload58_A clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_299_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19129_ net1184 _00170_ _00800_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[174\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13309__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout119_A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_329_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14506__B1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_342_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16322__A _06571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_239_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12532__A2 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_206_Left_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout390_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16041__B net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10543__B2 game.CPU.applesa.ab.absxs.body_x\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_318_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16976__B _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19515__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14285__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09715_ net1148 _03316_ game.CPU.applesa.ab.absxs.body_y\[20\] net895 _03956_ vssd1
+ vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__a221o_1
XANTENNA__15880__B net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11185__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12996__S net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout655_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_260_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout276_X net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18249__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17223__A2 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ net915 game.CPU.applesa.ab.check_walls.above.walls\[153\] game.CPU.applesa.ab.check_walls.above.walls\[157\]
+ net898 vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14037__A2 game.CPU.applesa.ab.check_walls.above.walls\[113\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_328_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_182_Right_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09577_ net1133 net820 vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__xor2_1
XFILLER_0_328_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16982__A1 _02462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19665__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12297__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_X net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_215_Left_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15104__C net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18980__Q game.CPU.applesa.ab.check_walls.above.walls\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20041__1365 vssd1 vssd1 vccd1 vccd1 _20041__1365/HI net1365 sky130_fd_sc_hd__conb_1
XFILLER_0_147_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16734__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13620__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11470_ net827 net261 _05349_ _05358_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10421_ _04192_ _04563_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__nor2_1
XFILLER_0_324_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_213_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14017__A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ net286 _07013_ net241 vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_189_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09893__X _04136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10352_ _00290_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__inv_2
XANTENNA__19045__CLK net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16503__Y _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13071_ game.writer.tracker.frame\[194\] game.writer.tracker.frame\[195\] net1030
+ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_224_Left_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10283_ net1458 _04473_ _04474_ game.CPU.applesa.ab.start_enable vssd1 vssd1 vccd1
+ vccd1 _01319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_264_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout91_X net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16232__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_295_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_292_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12022_ net820 net296 net290 net821 vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__a22o_1
XANTENNA__09924__B1 _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13720__B2 game.writer.tracker.frame\[200\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11376__A game.CPU.applesa.ab.check_walls.above.walls\[178\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16830_ net173 _02524_ net188 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__and3b_1
XFILLER_0_228_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14276__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 _04444_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_4
Xfanout581 net591 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11095__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout592 net595 vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_4
XANTENNA__15790__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16761_ net166 _02415_ net109 _02588_ net1621 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[182\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__13484__A0 _07048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13973_ _07844_ _07846_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_224_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18500_ net586 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__inv_2
X_12924_ _06697_ _06699_ net678 vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__mux2_1
XANTENNA__17214__A2 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15712_ _03289_ net344 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__xnor2_1
X_19480_ clknet_leaf_18_clk game.writer.tracker.next_frame\[75\] net1308 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[75\] sky130_fd_sc_hd__dfrtp_1
X_16692_ _02467_ net61 _02564_ net1576 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[138\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_220_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16422__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_244_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18431_ net601 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__inv_2
XFILLER_0_347_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12855_ game.writer.tracker.frame\[304\] game.writer.tracker.frame\[305\] net988
+ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__mux2_2
XANTENNA__11823__B _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15643_ net811 net437 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_233_Left_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15776__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11806_ net570 _05569_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__xnor2_1
X_15574_ game.CPU.kyle.L1.cnt_500hz\[9\] game.CPU.kyle.L1.cnt_500hz\[10\] game.CPU.kyle.L1.cnt_500hz\[11\]
+ _01586_ game.CPU.kyle.L1.cnt_500hz\[12\] vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__a41o_1
X_18362_ net596 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__inv_2
X_12786_ game.writer.tracker.frame\[346\] game.writer.tracker.frame\[347\] net1018
+ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12000__A game.CPU.applesa.ab.check_walls.above.walls\[165\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17313_ net176 _02409_ _02760_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[563\]
+ sky130_fd_sc_hd__a21o_1
X_14525_ _07398_ _07399_ _08370_ vssd1 vssd1 vccd1 vccd1 _08399_ sky130_fd_sc_hd__nand3_1
XFILLER_0_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11737_ game.CPU.applesa.ab.check_walls.above.walls\[108\] net392 _05618_ _05621_
+ _05624_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__o2111a_1
XANTENNA__19588__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18293_ net641 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
XANTENNA__16725__B2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16407__A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13530__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_313_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17244_ _02240_ _02257_ _02357_ net725 vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__o31a_1
X_14456_ game.CPU.applesa.ab.absxs.body_x\[15\] net1050 vssd1 vssd1 vccd1 vccd1 _08330_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_289_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11668_ net566 _05551_ _05555_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__o21ai_1
X_13407_ _06868_ _06878_ net680 vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17175_ _02472_ net73 _02724_ net1823 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[461\]
+ sky130_fd_sc_hd__a22o_1
X_10619_ net562 _04677_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__nand2_1
XANTENNA__15030__B net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10455__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14387_ game.CPU.applesa.ab.absxs.body_y\[6\] net951 vssd1 vssd1 vccd1 vccd1 _08261_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11599_ net800 net259 _05474_ _05475_ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16126_ _03466_ net346 net343 _03467_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_330_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13338_ _06601_ _06629_ net695 vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__mux2_1
XANTENNA__17150__A1 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_268_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15965__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10174__B game.CPU.applesa.ab.apple_possible\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16413__Y _02382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16057_ net1266 net474 net460 net1265 _02063_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__o221a_1
X_13269_ net209 _07134_ net284 vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_295_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13172__C1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19538__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15008_ net1220 net1248 net824 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__and3_1
XANTENNA__12514__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire456_A _08425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_284_Right_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19816_ clknet_leaf_37_clk game.writer.tracker.next_frame\[411\] net1349 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[411\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15981__A game.CPU.applesa.ab.check_walls.above.walls\[64\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_324_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_263_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_162_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19747_ clknet_leaf_24_clk game.writer.tracker.next_frame\[342\] net1340 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[342\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16959_ net168 net69 net94 _02658_ net1571 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[311\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__18562__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19688__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18069__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ _03738_ _03739_ _03741_ _03742_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__a211o_1
XANTENNA__17205__A2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19678_ clknet_leaf_34_clk game.writer.tracker.next_frame\[273\] net1319 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[273\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12829__B net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ net892 net799 _03443_ net1128 _03673_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_88_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18629_ clknet_leaf_16_clk _01046_ _00366_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_176_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16964__A1 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15767__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09362_ net1137 game.CPU.applesa.ab.check_walls.above.walls\[198\] vssd1 vssd1 vccd1
+ vccd1 _03605_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_43_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11789__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_353_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15519__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ net1091 game.CPU.applesa.ab.check_walls.above.walls\[82\] vssd1 vssd1 vccd1
+ vccd1 _03536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_11 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13440__S net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _06783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_33 _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_44 clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19068__CLK net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16036__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_306_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_278_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1145_A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13950__A1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13950__B2 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17141__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12580__A game.CPU.applesa.ab.absxs.body_x\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_274_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_273_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_262_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_251_Right_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10812__B _04702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19136__Q game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__A1 net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18905__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__B2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1100_X net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16241__A_N _06607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18975__Q game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ _03294_ net542 vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__nand2_1
XFILLER_0_329_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11643__B net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ net1109 game.CPU.applesa.ab.absxs.body_x\[16\] vssd1 vssd1 vccd1 vccd1 _03872_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_356_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16955__A1 _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12640_ game.CPU.applesa.ab.absxs.body_x\[17\] net377 game.CPU.applesa.twoapples.absxs.next_head\[3\]
+ _03282_ _06516_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__a221o_1
XFILLER_0_356_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_273_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_316_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12977__C1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12571_ game.CPU.applesa.ab.absxs.body_x\[17\] net377 net371 game.CPU.applesa.ab.absxs.body_x\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__o22a_1
XANTENNA__16707__A1 _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16227__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_195_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14310_ _08181_ _08182_ _08183_ vssd1 vssd1 vccd1 vccd1 _08184_ sky130_fd_sc_hd__or3_2
XFILLER_0_92_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11522_ net745 _05410_ _05409_ net568 vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__a2bb2o_1
X_15290_ game.CPU.applesa.twomode.counter_normal game.CPU.applesa.twomode.number\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08840_ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_324_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12474__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13616__S1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ game.CPU.applesa.ab.absxs.body_y\[113\] net865 net858 game.CPU.applesa.ab.absxs.body_y\[115\]
+ vssd1 vssd1 vccd1 vccd1 _08115_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_351_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11453_ game.CPU.applesa.ab.check_walls.above.walls\[78\] net257 net316 net813 vssd1
+ vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_190_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16514__X _02456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18442__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_312_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10404_ game.CPU.randy.f1.state\[3\] _04552_ _04550_ vssd1 vssd1 vccd1 vccd1 _01243_
+ sky130_fd_sc_hd__o21a_1
X_14172_ game.CPU.applesa.ab.absxs.body_x\[106\] net1056 vssd1 vssd1 vccd1 vccd1 _08046_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_296_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17132__A1 _02310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11384_ net784 net251 net318 game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1
+ vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__15785__B net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13123_ _06993_ _06995_ net696 vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__mux2_1
X_10335_ net1796 _04509_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__xnor2_1
X_18980_ net1201 _00205_ _00651_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14497__A2 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_284_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _06924_ _06926_ net687 vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__mux2_1
X_17931_ net659 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__inv_2
X_10266_ _04458_ _04377_ _04376_ _04401_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_237_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_226_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18585__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11704__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1310 net1314 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__clkbuf_4
X_12005_ net786 net294 net289 net787 vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__o22ai_1
XANTENNA__09373__A1 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1321 net1322 vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__clkbuf_4
XANTENNA__19830__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09373__B2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1332 net1333 vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__clkbuf_4
X_17862_ game.writer.updater.commands.count\[12\] game.writer.updater.commands.count\[13\]
+ _03178_ game.writer.updater.commands.count\[14\] vssd1 vssd1 vccd1 vccd1 _03183_
+ sky130_fd_sc_hd__a31o_1
Xfanout1343 net1348 vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__clkbuf_4
X_10197_ _04386_ _04388_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__nand2_1
XANTENNA__15009__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19601_ clknet_leaf_22_clk game.writer.tracker.next_frame\[196\] net1343 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[196\] sky130_fd_sc_hd__dfrtp_1
Xfanout1354 net1357 vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16643__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16813_ _02502_ net105 _02604_ net1788 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[219\]
+ sky130_fd_sc_hd__a22o_1
X_17793_ _03135_ net888 _03134_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__mux2_1
XANTENNA__15997__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19532_ clknet_leaf_23_clk game.writer.tracker.next_frame\[127\] net1344 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[127\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11834__A game.CPU.applesa.ab.check_walls.above.walls\[151\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_241_Left_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16744_ _02299_ net163 net101 _02583_ net1471 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[171\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_205_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_198_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13956_ net886 game.CPU.applesa.ab.check_walls.above.walls\[128\] game.CPU.applesa.ab.check_walls.above.walls\[129\]
+ net881 _07823_ vssd1 vssd1 vccd1 vccd1 _07830_ sky130_fd_sc_hd__a221o_1
XANTENNA_output32_A net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19463_ clknet_leaf_40_clk game.writer.tracker.next_frame\[58\] net1358 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[58\] sky130_fd_sc_hd__dfrtp_1
X_12907_ game.writer.tracker.frame\[50\] game.writer.tracker.frame\[51\] net1024 vssd1
+ vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__mux2_1
XANTENNA__11553__B net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15025__B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16675_ _02555_ _02556_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__and2_1
XANTENNA__16946__A1 _02390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13887_ net987 game.CPU.applesa.ab.check_walls.above.walls\[100\] vssd1 vssd1 vccd1
+ vccd1 _07761_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_319_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18414_ net626 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12838_ game.writer.tracker.frame\[318\] game.writer.tracker.frame\[319\] net1032
+ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_295_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15626_ game.CPU.applesa.ab.check_walls.above.walls\[187\] net457 vssd1 vssd1 vccd1
+ vccd1 _01638_ sky130_fd_sc_hd__xnor2_1
X_19394_ clknet_leaf_55_clk net1403 net1280 vssd1 vssd1 vccd1 vccd1 game.writer.control.detect4.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_347_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10169__B game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_237_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14421__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_335_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18345_ net593 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__inv_2
X_12769_ game.writer.tracker.frame\[114\] game.writer.tracker.frame\[115\] net1015
+ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__mux2_1
X_15557_ _01540_ _01575_ _01576_ _01470_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12665__A _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_334_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14508_ game.CPU.apple_location2\[3\] net1044 vssd1 vssd1 vccd1 vccd1 _08382_ sky130_fd_sc_hd__xor2_1
X_15488_ _01485_ _01488_ _01502_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18276_ net622 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_315_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12384__B net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_353_Right_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17227_ _02410_ net123 net121 _02737_ net1520 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[500\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_20_clk_X clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_342_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14439_ game.CPU.applesa.ab.absxs.body_y\[91\] net939 vssd1 vssd1 vccd1 vccd1 _08313_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_140_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16424__X _02390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14880__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13393__C1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_303_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19360__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09974__A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17123__A1 _02375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17158_ _02237_ net122 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__and2_1
XANTENNA__15695__B net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_326_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16109_ _02031_ _02034_ _02119_ _02120_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__or4b_1
XANTENNA__18928__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17089_ _02482_ net57 _02698_ game.writer.tracker.frame\[401\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[401\] sky130_fd_sc_hd__a22o_1
X_09980_ net1158 net848 _04206_ vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_228_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10913__A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_35_clk_X clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_248_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10632__B net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14104__B game.CPU.applesa.ab.check_walls.above.walls\[53\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_139_Left_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13791__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_271_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20040__1364 vssd1 vssd1 vccd1 vccd1 _20040__1364/HI net1364 sky130_fd_sc_hd__conb_1
XANTENNA__13435__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout186_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_329_Left_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13999__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13999__B2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_337_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09414_ net1128 game.CPU.applesa.ab.absxs.body_y\[99\] vssd1 vssd1 vccd1 vccd1 _03657_
+ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout1095_A game.CPU.applesa.ab.snake_head_x\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_90_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ net1142 game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1 _03588_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout520_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__A1 game.CPU.applesa.ab.absxs.body_y\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout141_X net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout239_X net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09276_ game.CPU.walls.rand_wall.count_luck\[0\] vssd1 vssd1 vccd1 vccd1 _03523_
+ sky130_fd_sc_hd__inv_2
XANTENNA__19703__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_340_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_320_Right_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15886__A game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_338_Left_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_306_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1050_X net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18262__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1148_X net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13923__A1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13923__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_348_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16607__A_N _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_210_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10737__A1 game.CPU.applesa.ab.absxs.body_y\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_160_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout987_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10737__B2 game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19853__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14479__A2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout99_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ game.CPU.applesa.enable_in game.CPU.applesa.twoapples.x_final\[0\] _03212_
+ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_356_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10051_ game.CPU.applesa.twoapples.count_luck\[7\] game.CPU.applesa.twoapples.count_luck\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__or2_1
XANTENNA__13782__S0 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16510__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_356_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13810_ _07682_ _07683_ net497 vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_242_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_242_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14790_ net1754 _08604_ _08607_ vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_215_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09658__A2 game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_221_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13741_ game.writer.tracker.frame\[241\] game.writer.tracker.frame\[243\] game.writer.tracker.frame\[244\]
+ game.writer.tracker.frame\[242\] net978 net1027 vssd1 vssd1 vccd1 vccd1 _07615_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09124__A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10953_ _04832_ _04833_ _04835_ _04836_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a22o_1
XANTENNA__16928__A1 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17050__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16460_ net1883 _02414_ _02416_ net137 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[54\]
+ sky130_fd_sc_hd__a22o_1
X_13672_ game.writer.tracker.frame\[461\] game.writer.tracker.frame\[463\] game.writer.tracker.frame\[464\]
+ game.writer.tracker.frame\[462\] net974 net1010 vssd1 vssd1 vccd1 vccd1 _07546_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_195_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10884_ _04779_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__or2_1
XANTENNA__14403__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15600__A1 game.CPU.applesa.ab.check_walls.above.walls\[113\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13837__S1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_317_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15411_ _08901_ _01437_ _01438_ _08934_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__o211a_1
XFILLER_0_210_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ _06303_ _06305_ _06312_ _06498_ _06499_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__o311a_1
X_16391_ _02274_ _02365_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__or2_1
XFILLER_0_183_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_316_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09778__B game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_23_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_241_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15342_ game.writer.updater.commands.cmd_num\[1\] _03366_ _08882_ _08883_ vssd1 vssd1
+ vccd1 vccd1 _08884_ sky130_fd_sc_hd__o31a_1
X_18130_ net578 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__inv_2
X_12554_ game.CPU.applesa.ab.absxs.body_x\[86\] net370 net528 game.CPU.applesa.ab.absxs.body_x\[87\]
+ _06430_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__o221a_1
XFILLER_0_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19383__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_310_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13868__X _07742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11505_ net785 net250 _05392_ _05393_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__a211oi_1
X_15273_ _08827_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__inv_2
X_18061_ net613 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__inv_2
X_12485_ _06353_ _06355_ _06361_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__or3b_1
XFILLER_0_108_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16244__X _02252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17012_ _02499_ net90 net558 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_232_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14224_ game.CPU.applesa.ab.absxs.body_x\[42\] net1059 vssd1 vssd1 vccd1 vccd1 _08098_
+ sky130_fd_sc_hd__nand2_1
X_11436_ net567 _05319_ _05320_ _05324_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__a211oi_1
XANTENNA__17105__A1 _02574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10728__A1 game.CPU.applesa.ab.absxs.body_y\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_123_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16404__B net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14155_ net1161 net993 vssd1 vssd1 vccd1 vccd1 _08029_ sky130_fd_sc_hd__xor2_1
XFILLER_0_104_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11367_ net745 _05255_ _05253_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__a21o_1
XFILLER_0_238_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13106_ net508 _06979_ _06978_ net210 vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__o211a_1
XFILLER_0_237_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10318_ _04487_ _04496_ _04499_ net739 net2030 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__a32o_1
X_18963_ net1199 _00276_ _00634_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_14086_ net1059 game.CPU.applesa.ab.check_walls.above.walls\[90\] vssd1 vssd1 vccd1
+ vccd1 _07960_ sky130_fd_sc_hd__xor2_1
XANTENNA__13678__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11298_ _05141_ _05142_ _05187_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__or3_1
X_13037_ net484 _06908_ _06910_ net275 vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__a211o_1
XFILLER_0_266_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17914_ net605 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__inv_2
X_10249_ net774 net770 vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__nand2_2
X_18894_ clknet_leaf_2_clk _01266_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1140 net1143 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_266_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1151 net1152 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_321_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17845_ net182 _03168_ game.writer.updater.commands.count\[9\] vssd1 vssd1 vccd1
+ vccd1 _03171_ sky130_fd_sc_hd__o21bai_1
Xfanout1162 game.CPU.applesa.twoapples.logic_enable vssd1 vssd1 vccd1 vccd1 net1162
+ sky130_fd_sc_hd__buf_2
Xfanout1173 net1174 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__clkbuf_2
Xfanout1184 net1190 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__buf_2
Xfanout1195 game.CPU.walls.rand_wall.good_spot vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__buf_2
X_17776_ _03125_ _03126_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14988_ net1227 net1254 game.CPU.applesa.ab.check_walls.above.walls\[16\] vssd1 vssd1
+ vccd1 vccd1 _00204_ sky130_fd_sc_hd__and3_1
X_19515_ clknet_leaf_14_clk game.writer.tracker.next_frame\[110\] net1283 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[110\] sky130_fd_sc_hd__dfrtp_1
X_16727_ net161 _02434_ net106 _02578_ net1642 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[159\]
+ sky130_fd_sc_hd__a32o_1
X_13939_ net1065 game.CPU.applesa.ab.check_walls.above.walls\[65\] vssd1 vssd1 vccd1
+ vccd1 _07813_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_18_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11456__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16419__X _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_240_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_62_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_338_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19446_ clknet_leaf_47_clk game.writer.tracker.next_frame\[41\] net1298 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[41\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09969__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16658_ net153 net128 _02422_ _02546_ net1782 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[121\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__18600__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19726__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15609_ game.CPU.applesa.ab.absxs.body_y\[33\] net340 vssd1 vssd1 vccd1 vccd1 _01621_
+ sky130_fd_sc_hd__nand2_1
X_19377_ clknet_leaf_3_clk _01383_ _00958_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.snake_head_y\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_16589_ net1849 _02505_ _02506_ net126 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[93\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ net832 vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__inv_2
X_18328_ net616 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_157_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_332_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_322_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14158__A1 net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_170_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09061_ game.CPU.applesa.ab.absxs.body_y\[45\] vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__inv_2
XANTENNA__19876__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_288_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10119__S _04311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18259_ net622 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XANTENNA__18750__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_301_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload40_A clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 game.writer.tracker.frame\[19\] vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10719__A1 game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_330_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold612 game.writer.tracker.frame\[29\] vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap331 _08451_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11739__A game.CPU.applesa.ab.check_walls.above.walls\[157\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold623 game.CPU.kyle.L1.currentState\[2\] vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13381__A2 _07241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold634 game.writer.tracker.frame\[555\] vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout101_A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold645 game.CPU.randy.f1.a1.count\[14\] vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 game.writer.tracker.frame\[9\] vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14115__A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_147_Left_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold667 game.writer.tracker.frame\[242\] vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13118__C1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16855__B1 _02623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09209__A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09963_ net903 _04190_ _04192_ _04191_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__a31o_1
XANTENNA__11458__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16601__Y _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13954__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17426__A _02779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16870__A3 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09894_ _03584_ _03587_ _04130_ _04132_ _04136_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__o2111a_1
XANTENNA__16330__A _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_168_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__C net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_181_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17280__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_X net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14488__C _08358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_A _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12289__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12644__A1 _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13841__B1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout735_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_X net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18257__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_156_Left_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1098_X net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_257_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_270_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout902_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1265_X net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_346_Left_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09328_ _03568_ _03570_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__nand2_1
XANTENNA__15112__C game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11080__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ game.CPU.randy.counter1.count\[6\] vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_334_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12270_ game.CPU.applesa.ab.check_walls.above.walls\[111\] net423 vssd1 vssd1 vccd1
+ vccd1 _06156_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout892_X net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_165_Left_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17099__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09576__A1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ game.CPU.applesa.ab.absxs.body_y\[39\] net400 vssd1 vssd1 vccd1 vccd1 _05111_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09576__B2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11649__A game.CPU.applesa.ab.check_walls.above.walls\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14025__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11383__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13109__C1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_268_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_287_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16846__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09119__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ game.CPU.applesa.ab.absxs.body_x\[98\] net411 net400 game.CPU.applesa.ab.absxs.body_y\[99\]
+ _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__o221a_1
XANTENNA__11368__B net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_281_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16511__Y _02454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10103_ _04252_ _04258_ _04310_ _04256_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.good_spot_next
+ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_355_Left_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13755__S0 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15960_ _03395_ game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 _01972_ sky130_fd_sc_hd__nor2_1
X_11083_ _04969_ _04972_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__nand2_1
XANTENNA__16861__A3 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14911_ net1174 _08430_ _08687_ vssd1 vssd1 vccd1 vccd1 _08688_ sky130_fd_sc_hd__a21oi_1
X_10034_ _04217_ _04223_ _04231_ _04241_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__or4_1
XANTENNA__12883__A1 game.writer.tracker.frame\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15891_ _01895_ _01896_ _01897_ _01902_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__or4_2
X_17630_ game.CPU.kyle.L1.cnt_20ms\[16\] game.CPU.kyle.L1.cnt_20ms\[15\] _03032_ vssd1
+ vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__and3_1
XANTENNA__09125__Y _03374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14842_ _04332_ _08639_ _08640_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[5\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_236_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18623__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14085__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19749__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_174_Left_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_349_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17561_ net1461 _08808_ _02986_ net429 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14773_ _08584_ _08586_ _08592_ _08593_ vssd1 vssd1 vccd1 vccd1 _08594_ sky130_fd_sc_hd__o31a_1
X_11985_ _05267_ _05268_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__nand2_1
XANTENNA__13832__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19300_ clknet_leaf_56_clk game.CPU.applesa.ab.check_walls.collision_leftn _00915_
+ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.collision_left sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16512_ net149 net128 _02454_ _02446_ net1800 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[68\]
+ sky130_fd_sc_hd__a32o_1
X_13724_ net492 _07596_ _07597_ vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__and3_1
X_10936_ _03356_ net404 vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_15_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17492_ net1258 net1259 game.CPU.speed1.Qa\[0\] net427 vssd1 vssd1 vccd1 vccd1 _02921_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_156_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_357_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_317_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_292_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19231_ clknet_leaf_57_clk net1418 _00869_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.normal1.number\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_16443_ net171 _02403_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__nor2_4
XFILLER_0_156_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19899__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13655_ game.writer.tracker.frame\[1\] game.writer.tracker.frame\[3\] game.writer.tracker.frame\[4\]
+ game.writer.tracker.frame\[2\] net969 net1002 vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__mux4_1
X_10867_ _03516_ game.CPU.randy.counter1.count1\[1\] _04762_ vssd1 vssd1 vccd1 vccd1
+ _04770_ sky130_fd_sc_hd__a21o_1
XANTENNA__18773__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14388__B2 game.CPU.applesa.ab.absxs.body_y\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_234_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12606_ game.CPU.applesa.ab.absxs.body_y\[62\] net521 net361 game.CPU.applesa.ab.absxs.body_y\[60\]
+ _06376_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__o221a_1
X_19162_ clknet_leaf_67_clk _01282_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count_luck\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_13586_ game.writer.tracker.frame\[341\] game.writer.tracker.frame\[343\] game.writer.tracker.frame\[344\]
+ game.writer.tracker.frame\[342\] net979 net1029 vssd1 vssd1 vccd1 vccd1 _07460_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__17326__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16374_ _02284_ _02313_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__nand2_2
XANTENNA__15022__C game.CPU.applesa.ab.check_walls.above.walls\[50\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10798_ game.CPU.applesa.ab.absxs.body_y\[35\] _04696_ _04697_ game.CPU.applesa.ab.absxs.body_y\[31\]
+ vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_304_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10949__B2 game.CPU.applesa.ab.absxs.body_y\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18113_ net583 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_313_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15325_ game.CPU.applesa.twomode.number\[6\] _08864_ vssd1 vssd1 vccd1 vccd1 _08869_
+ sky130_fd_sc_hd__and2_1
X_12537_ game.CPU.applesa.ab.absxs.body_x\[43\] net531 vssd1 vssd1 vccd1 vccd1 _06414_
+ sky130_fd_sc_hd__xnor2_1
X_19093_ net1178 _00130_ _00764_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[138\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_297_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19129__CLK net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_183_Left_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18044_ net659 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__inv_2
X_12468_ game.CPU.applesa.ab.absxs.body_y\[12\] net361 vssd1 vssd1 vccd1 vccd1 _06345_
+ sky130_fd_sc_hd__xnor2_1
X_15256_ _08813_ _01264_ vssd1 vssd1 vccd1 vccd1 _08814_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09567__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14207_ _08073_ _08074_ _08079_ _08080_ vssd1 vssd1 vccd1 vccd1 _08081_ sky130_fd_sc_hd__or4_1
XANTENNA__09567__B2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11419_ net566 _05301_ _05303_ _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__a211o_1
X_15187_ _08760_ game.CPU.walls.enable_in2 vssd1 vssd1 vccd1 vccd1 _08762_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12007__X _05894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12399_ game.CPU.applesa.ab.absxs.body_y\[95\] net364 vssd1 vssd1 vccd1 vccd1 _06276_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__11382__A1_N net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11374__A1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12571__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14138_ net1061 _03402_ _03403_ net963 vssd1 vssd1 vccd1 vccd1 _08012_ sky130_fd_sc_hd__a22o_1
XFILLER_0_238_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15973__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16301__A2 _02300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19995_ clknet_leaf_44_clk _01419_ net1304 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10182__B game.CPU.applesa.ab.apple_possible\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19279__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_245_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09319__A1 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_288_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14069_ net1075 _03378_ _03380_ net956 _07942_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18946_ net1175 _00075_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.counter sky130_fd_sc_hd__dfxtp_2
XFILLER_0_225_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_3_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__12323__B1 _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18877_ clknet_leaf_5_clk game.CPU.randy.f1.c1.innerCount\[7\] _00572_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10910__B game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_192_Left_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17828_ _03158_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__inv_2
XFILLER_0_206_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14076__B1 game.CPU.applesa.ab.YMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17759_ game.CPU.applesa.twoapples.count_luck\[2\] _03113_ game.CPU.applesa.twoapples.count_luck\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_334_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09699__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19429_ clknet_leaf_41_clk game.writer.tracker.next_frame\[24\] net1332 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10638__A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout149_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17317__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09113_ net1272 vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13949__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16325__A net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout316_A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14580__B1_N net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ game.CPU.applesa.ab.absxs.body_y\[102\] vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12572__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold420 game.writer.tracker.frame\[345\] vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_345_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout104_X net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold431 game.CPU.randy.f1.c1.count\[12\] vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_276_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold442 game.writer.tracker.frame\[423\] vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1225_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold453 game.writer.tracker.frame\[41\] vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 game.writer.tracker.frame\[93\] vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11188__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold475 game.CPU.kyle.L1.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold486 game.CPU.kyle.L1.currentState\[1\] vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout685_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_8
Xhold497 game.writer.tracker.frame\[59\] vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 net913 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__buf_2
XANTENNA__14303__A1 game.CPU.applesa.ab.absxs.body_y\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13737__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_284_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout922 net923 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_4
XANTENNA__16843__A3 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09946_ net1116 _04178_ net1115 vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout1013_X net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout933 net934 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__buf_2
XANTENNA__18646__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout944 net945 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14499__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12314__B1 _06150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout955 net956 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_2
Xfanout966 net973 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__clkbuf_2
Xfanout977 net982 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_232_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ _03711_ _03716_ _04118_ _04119_ _03638_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout852_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16995__A _02455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout988 net989 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16056__A1 net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout999 net1000 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09730__A1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16056__B2 net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09730__B2 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19454__RESET_B net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15107__C game.CPU.applesa.ab.check_walls.above.walls\[135\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10340__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18983__Q game.CPU.applesa.ab.check_walls.above.walls\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12617__A1 net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18796__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__A2_N net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11932__A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11770_ _03450_ net299 vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17556__A1 _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11651__B net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10721_ game.CPU.applesa.ab.absxs.body_y\[45\] _04640_ _04641_ game.CPU.applesa.ab.absxs.body_y\[41\]
+ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_354_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10548__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13440_ _06925_ _06935_ net687 vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__mux2_1
XANTENNA__09896__X _04139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10652_ _04585_ _04607_ _04156_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__o21ai_4
XANTENNA__10267__B net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09797__A1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13371_ _07243_ _07244_ net501 vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__mux2_1
XANTENNA__09797__B2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10583_ game.CPU.applesa.ab.absxs.body_x\[114\] _04663_ _04664_ game.CPU.applesa.ab.absxs.body_x\[110\]
+ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__a22o_1
XANTENNA__16235__A _02238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15110_ net1204 net1231 game.CPU.applesa.ab.check_walls.above.walls\[138\] vssd1
+ vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12322_ _06204_ _06205_ _06206_ _06207_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.collision
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_152_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16090_ _02092_ _02101_ _02093_ _02097_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__or4b_2
XANTENNA__16531__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_279_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09549__A1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11379__A game.CPU.applesa.ab.check_walls.above.walls\[177\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15041_ net1219 net1248 net815 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__and3_1
XANTENNA__19421__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09549__B2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ _05980_ _05981_ _06137_ _06138_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__or4_1
XFILLER_0_133_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11204_ game.CPU.applesa.ab.absxs.body_x\[92\] net326 vssd1 vssd1 vccd1 vccd1 _05094_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__11098__B net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12184_ game.CPU.applesa.ab.check_walls.above.walls\[62\] net419 vssd1 vssd1 vccd1
+ vccd1 _06070_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15793__B net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20044__X net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16295__A1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18800_ clknet_leaf_71_clk game.CPU.clock1.next_counter\[3\] _00537_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13728__S0 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ game.CPU.applesa.ab.absxs.body_x\[68\] net325 vssd1 vssd1 vccd1 vccd1 _05025_
+ sky130_fd_sc_hd__nand2_1
X_19780_ clknet_leaf_24_clk game.writer.tracker.next_frame\[375\] net1344 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[375\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_208_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10570__X _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__B game.CPU.applesa.ab.absxs.body_x\[40\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16992_ _02475_ net88 _02668_ net1799 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[334\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13502__C1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19571__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_196_Right_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18731_ clknet_leaf_13_clk _01148_ _00468_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[113\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11826__B net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066_ _03279_ net319 vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__nor2_1
X_15943_ net820 net432 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__nor2_1
XANTENNA__14202__B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13881__X _07755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17244__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ net1081 _04224_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__and2_1
XANTENNA__09721__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09721__B2 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18662_ clknet_leaf_64_clk _01079_ _00399_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[84\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15874_ _03278_ net343 net444 game.CPU.applesa.ab.absxs.body_y\[25\] vssd1 vssd1
+ vccd1 vccd1 _01886_ sky130_fd_sc_hd__a22o_1
XANTENNA__17795__B2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17613_ _03023_ _03024_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_240_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ game.CPU.randy.counter1.count\[17\] _08628_ vssd1 vssd1 vccd1 vccd1 _08630_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_263_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18593_ clknet_leaf_50_clk _01013_ _00330_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[66\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_230_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17544_ _02948_ _02966_ _02969_ _02970_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__or4_1
X_14756_ net54 _08577_ _08578_ vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__and3_1
X_11968_ game.CPU.applesa.ab.check_walls.above.walls\[148\] net551 vssd1 vssd1 vccd1
+ vccd1 _05855_ sky130_fd_sc_hd__nand2_1
XANTENNA__09312__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_317_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13707_ net226 _07576_ _07580_ net277 vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__o211a_1
XANTENNA__15033__B net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11292__B1 _05181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_345_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10919_ net1166 _04391_ _04813_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__a21o_1
X_17475_ _02898_ _02900_ _02903_ _02893_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__a22o_1
X_11899_ net751 _05410_ _05415_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__o21ai_1
X_14687_ _04347_ _08491_ game.CPU.randy.counter1.count1\[14\] vssd1 vssd1 vccd1 vccd1
+ _08526_ sky130_fd_sc_hd__a21o_1
X_19214_ net1168 _00026_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_possible\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_16426_ net219 _02310_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__and2_2
XFILLER_0_144_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13638_ _07510_ _07511_ net495 vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__mux2_1
XANTENNA__15968__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_305_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13769__A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19145_ net1188 _00188_ _00816_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[190\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13584__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16357_ net136 _02258_ _02341_ _02338_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[26\]
+ sky130_fd_sc_hd__a31o_1
X_13569_ game.writer.tracker.frame\[333\] game.writer.tracker.frame\[335\] game.writer.tracker.frame\[336\]
+ game.writer.tracker.frame\[334\] net968 net999 vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_313_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15308_ game.CPU.applesa.twomode.number\[3\] _08849_ vssd1 vssd1 vccd1 vccd1 _08855_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19076_ net1179 _00112_ _00747_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[121\]
+ sky130_fd_sc_hd__dfrtp_4
X_16288_ net479 net836 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__nand2_1
XANTENNA__15984__A game.CPU.applesa.ab.check_walls.above.walls\[65\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_18027_ net647 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__inv_2
XFILLER_0_301_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15239_ game.CPU.kyle.L1.cnt_500hz\[0\] game.CPU.kyle.L1.cnt_500hz\[1\] vssd1 vssd1
+ vccd1 vccd1 _08800_ sky130_fd_sc_hd__nand2_1
XANTENNA__16432__X _02395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_288_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18669__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19914__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19965__RESET_B net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout207 net208 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_2
X_09800_ net1083 _03437_ net800 net907 vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__a22o_1
XANTENNA__09960__A1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_238_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout218 _06592_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_4
Xfanout229 net232 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_2
X_19978_ clknet_leaf_42_clk game.writer.tracker.next_frame\[573\] net1326 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[573\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14297__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11736__B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09731_ net1091 _03275_ _03276_ net1098 vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__a22o_1
X_18929_ clknet_leaf_5_clk net1411 _00613_ vssd1 vssd1 vccd1 vccd1 game.CPU.right_button.eD1.D
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_340_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09712__A1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09712__B2 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ net1095 _03244_ _03313_ net1161 _03904_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__a221o_1
XFILLER_0_307_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09593_ net1133 game.CPU.applesa.ab.absxs.body_y\[75\] vssd1 vssd1 vccd1 vccd1 _03836_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__19341__D game.CPU.applesa.twoapples.absxs.collision vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17538__A1 net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16039__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11283__B1 _04930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_254_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout433_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16761__A2 _02415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_279_Left_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_176_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_351_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11035__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13679__A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19444__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout600_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1342_A net1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_X net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_298_Right_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ game.CPU.applesa.ab.absxs.body_x\[33\] vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1130_X net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18270__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1228_X net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19594__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 game.writer.tracker.frame\[107\] vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 game.writer.tracker.frame\[297\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_348_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_265_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 game.writer.tracker.frame\[488\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16502__B net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold283 game.writer.tracker.frame\[531\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 game.writer.tracker.frame\[378\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_207_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_348_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout81_A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14288__B1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout730 net738 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_288_Left_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_272_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout741 _04485_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_217_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09929_ net1100 net848 _04168_ vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11646__B net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout763 net764 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_129_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout774 net776 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_304_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout785 game.CPU.applesa.ab.check_walls.above.walls\[172\] vssd1 vssd1 vccd1 vccd1
+ net785 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09703__A1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout796 game.CPU.applesa.ab.check_walls.above.walls\[119\] vssd1 vssd1 vccd1 vccd1
+ net796 sky130_fd_sc_hd__clkbuf_4
X_20049_ net1368 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
X_12940_ _06741_ _06742_ net677 vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__mux2_1
XANTENNA__09703__B2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12871_ game.writer.tracker.frame\[36\] game.writer.tracker.frame\[37\] net1003 vssd1
+ vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__mux2_1
X_14610_ game.CPU.clock1.counter\[7\] game.CPU.clock1.counter\[8\] _08460_ vssd1 vssd1
+ vccd1 vccd1 _08464_ sky130_fd_sc_hd__and3_1
XANTENNA__15134__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11662__A game.CPU.applesa.ab.check_walls.above.walls\[123\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11822_ _05672_ _05679_ _05689_ _05699_ _05709_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_202_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _03398_ net345 net442 net822 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__a22o_1
XANTENNA__17529__B2 game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_276_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12477__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11381__B net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ net569 _05388_ _05639_ _05640_ _05382_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__o2111a_1
X_14541_ game.CPU.walls.rand_wall.logic_enable _04808_ vssd1 vssd1 vccd1 vccd1 _08413_
+ sky130_fd_sc_hd__nor2_2
XFILLER_0_28_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11813__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12494__A2_N net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_297_Left_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_218_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18445__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10704_ game.CPU.applesa.ab.absxs.body_y\[70\] _04625_ _04626_ game.CPU.applesa.ab.absxs.body_y\[66\]
+ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__a22o_1
X_17260_ net224 net136 _02619_ net722 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__o31a_1
XFILLER_0_354_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14472_ game.CPU.applesa.ab.absxs.body_y\[10\] net953 vssd1 vssd1 vccd1 vccd1 _08346_
+ sky130_fd_sc_hd__xnor2_1
X_11684_ net744 _05568_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__nor2_1
XANTENNA__15788__B net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_342_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12764__Y _06638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16752__A2 _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16211_ _01944_ _01947_ _01950_ _02222_ _01838_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__o311a_1
XANTENNA__13566__A2 game.writer.tracker.frame\[368\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13423_ _06986_ _06989_ _07001_ _06990_ net696 net482 vssd1 vssd1 vccd1 vccd1 _07297_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ net932 game.CPU.applesa.ab.absxs.body_x\[47\] net561 _04685_ vssd1 vssd1
+ vccd1 vccd1 _01118_ sky130_fd_sc_hd__a31o_1
XFILLER_0_165_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17191_ net149 _02498_ net78 _02728_ net1512 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[473\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_180_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11577__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13354_ _07226_ _07227_ net229 vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16142_ game.CPU.applesa.ab.absxs.body_y\[77\] net448 net432 game.CPU.applesa.ab.absxs.body_y\[79\]
+ _02153_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__o221a_1
XFILLER_0_141_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_265_Right_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10566_ game.CPU.applesa.ab.absxs.body_x\[13\] _04653_ _04654_ game.CPU.applesa.ab.absxs.body_x\[9\]
+ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19049__Q game.CPU.applesa.ab.check_walls.above.walls\[94\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12305_ net820 net423 vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__nor2_1
X_13285_ net209 _07158_ net277 vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__a21o_1
XANTENNA__12780__X _06654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16073_ game.CPU.applesa.ab.absxs.body_y\[84\] net449 vssd1 vssd1 vccd1 vccd1 _02085_
+ sky130_fd_sc_hd__xnor2_1
X_10497_ _03197_ _04578_ net1119 net1124 vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_307_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19901_ clknet_leaf_15_clk game.writer.tracker.next_frame\[496\] net1288 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[496\] sky130_fd_sc_hd__dfrtp_1
X_12236_ _06118_ _06121_ _06119_ _06120_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__or4b_2
X_15024_ net1222 net1250 game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1
+ vccd1 vccd1 _00244_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_287_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_258_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_310_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16412__B _02340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_229_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19832_ clknet_leaf_33_clk game.writer.tracker.next_frame\[427\] net1325 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[427\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18961__CLK net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12167_ game.CPU.applesa.ab.check_walls.above.walls\[157\] net386 vssd1 vssd1 vccd1
+ vccd1 _06054_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_258_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14279__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_242_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11118_ game.CPU.applesa.ab.absxs.body_x\[18\] net410 vssd1 vssd1 vccd1 vccd1 _05008_
+ sky130_fd_sc_hd__xnor2_1
X_19763_ clknet_leaf_30_clk game.writer.tracker.next_frame\[358\] net1292 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[358\] sky130_fd_sc_hd__dfrtp_1
X_16975_ net152 _02452_ net90 _02662_ net1639 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[323\]
+ sky130_fd_sc_hd__a32o_1
X_12098_ _05982_ _05983_ _05984_ _05977_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a31o_1
XANTENNA__15028__B net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_274_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18714_ clknet_leaf_64_clk _01131_ _00451_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[80\]
+ sky130_fd_sc_hd__dfrtp_4
X_11049_ game.CPU.applesa.ab.absxs.body_y\[80\] net533 vssd1 vssd1 vccd1 vccd1 _04939_
+ sky130_fd_sc_hd__xor2_1
X_15926_ _01929_ _01930_ _01935_ _01936_ _01937_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a221o_1
X_19694_ clknet_leaf_30_clk game.writer.tracker.next_frame\[289\] net1292 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[289\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_max_cap66_X net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11501__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19317__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 gpio_in[5] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_274_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18645_ clknet_leaf_53_clk _01062_ _00382_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[47\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15779__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15857_ _01862_ _01863_ _01864_ _01866_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_318_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14808_ game.CPU.randy.counter1.count\[11\] game.CPU.randy.counter1.count\[10\] _08616_
+ vssd1 vssd1 vccd1 vccd1 _08619_ sky130_fd_sc_hd__and3_1
X_18576_ clknet_leaf_65_clk _00996_ _00313_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[33\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_349_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15788_ game.CPU.applesa.ab.absxs.body_x\[74\] net469 vssd1 vssd1 vccd1 vccd1 _01800_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_160_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16991__A2 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12387__B net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09042__A game.CPU.applesa.ab.absxs.body_x\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17527_ _04482_ _02851_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11265__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19467__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15979__A game.CPU.applesa.ab.check_walls.above.walls\[66\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14739_ game.CPU.randy.counter1.count1\[12\] _08565_ vssd1 vssd1 vccd1 vccd1 _08567_
+ sky130_fd_sc_hd__and2_1
XANTENNA__14883__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_320_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09977__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17458_ _02770_ _02773_ _02775_ _02786_ _02813_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__o311a_1
XFILLER_0_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14203__B1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13557__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16409_ net1838 _02371_ _02378_ net115 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[41\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17389_ net1274 _02782_ net428 vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__and3_1
XFILLER_0_333_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19128_ net1183 _00169_ _00799_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[173\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_41_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09630__B1 game.CPU.applesa.ab.absxs.body_y\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_299_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_232_Right_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_286_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19059_ net1186 _00093_ _00730_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[104\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_329_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_285_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18090__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_342_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10922__Y game.CPU.applesa.ab.absxs.next_head\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_273_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16322__B net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Left_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09933__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_254_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11740__B2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11466__B net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17208__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_310_Left_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09714_ net1092 _03249_ _03250_ net1100 _03955_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__a221o_1
XFILLER_0_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_260_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09645_ net910 game.CPU.applesa.ab.check_walls.above.walls\[152\] game.CPU.applesa.ab.check_walls.above.walls\[154\]
+ net920 vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19422__Q game.writer.tracker.frame\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1292_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09576_ net892 game.CPU.applesa.ab.check_walls.above.walls\[44\] net821 net903 _03818_
+ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__a221o_1
XFILLER_0_334_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12297__B net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16982__A2 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10059__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13796__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1080_X net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16734__A2 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_350_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_324_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ game.CPU.left_button.eD1.Q2 game.CPU.left_button.eD1.Q1 _04153_ _04563_ vssd1
+ vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__and4b_1
XFILLER_0_190_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15120__C net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16498__A1 game.writer.tracker.frame\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_213_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11964__D1 _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11609__A2_N net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16498__B2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10351_ game.CPU.walls.rand_wall.counter2\[0\] _04517_ game.CPU.walls.rand_wall.counter2\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_189_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16513__A _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13070_ game.writer.tracker.frame\[196\] game.writer.tracker.frame\[197\] net1030
+ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_249_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10282_ net851 game.CPU.applesa.ab.y_final\[3\] game.CPU.applesa.ab.good_spot_next
+ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout972_X net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10832__Y _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12021_ net820 net296 net290 net821 vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_264_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09924__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13720__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14033__A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout84_X net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09127__A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11376__B net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 game.CPU.button_reset_in vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_4
Xfanout571 net572 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__buf_2
XANTENNA__13872__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16760_ net185 _02412_ net109 _02588_ net1640 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[181\]
+ sky130_fd_sc_hd__a32o_1
Xfanout582 net585 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_4
Xfanout593 net595 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_2
X_13972_ net887 game.CPU.applesa.ab.check_walls.above.walls\[80\] net808 net857 _07845_
+ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__o221a_1
XANTENNA__08966__A game.CPU.applesa.ab.absxs.body_y\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15711_ _03292_ net272 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__xnor2_1
X_12923_ net502 _06796_ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_224_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16691_ _02303_ _02561_ net719 vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__o21a_1
XANTENNA__16422__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11392__A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18430_ net586 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__inv_2
X_15642_ game.CPU.applesa.ab.check_walls.above.walls\[73\] net472 vssd1 vssd1 vccd1
+ vccd1 _01654_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_244_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12854_ _06724_ _06725_ _06727_ _06726_ net476 net677 vssd1 vssd1 vccd1 vccd1 _06728_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_213_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_334_Right_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18361_ net597 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11805_ net750 _05568_ _05572_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12775__X _06649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15573_ game.CPU.kyle.L1.cnt_500hz\[5\] game.CPU.kyle.L1.cnt_500hz\[6\] game.CPU.kyle.L1.cnt_500hz\[7\]
+ game.CPU.kyle.L1.cnt_500hz\[8\] vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__a31o_1
X_12785_ game.writer.tracker.frame\[348\] game.writer.tracker.frame\[349\] net1018
+ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__mux2_1
XANTENNA__12000__B net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17312_ _02276_ _02535_ game.writer.tracker.frame\[563\] net732 vssd1 vssd1 vccd1
+ vccd1 _02760_ sky130_fd_sc_hd__o211a_1
XFILLER_0_260_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14524_ _07164_ _07400_ _07742_ _08028_ vssd1 vssd1 vccd1 vccd1 _08398_ sky130_fd_sc_hd__or4_1
X_11736_ game.CPU.applesa.ab.check_walls.above.walls\[109\] net307 vssd1 vssd1 vccd1
+ vccd1 _05624_ sky130_fd_sc_hd__xor2_1
XANTENNA__16186__B1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18292_ net641 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16407__B _02376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17243_ _02553_ net79 _02741_ game.writer.tracker.frame\[512\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[512\] sky130_fd_sc_hd__a22o_1
XANTENNA__13539__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_313_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14455_ _08327_ _08328_ vssd1 vssd1 vccd1 vccd1 _08329_ sky130_fd_sc_hd__nand2_1
X_11667_ net742 _05552_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_289_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ net697 _06882_ _07279_ net484 vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17174_ _02471_ net74 _02724_ net1545 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[460\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10618_ _04631_ _04358_ _04600_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__or3b_1
X_11598_ net800 net259 _05486_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__o21ai_1
X_14386_ _03226_ net1072 net941 _03215_ vssd1 vssd1 vccd1 vccd1 _08260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_268_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_269_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16125_ _03464_ net269 net459 game.CPU.applesa.ab.check_walls.above.walls\[163\]
+ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a22o_1
X_13337_ _06628_ _06630_ net695 vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10549_ _03278_ net330 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17150__A2 _02693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19557__RESET_B net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16423__A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10773__A2 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11749__A1_N game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16056_ net1266 net472 net460 net1265 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__a22o_1
X_13268_ net694 _07141_ _07138_ net221 vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__o211a_1
XFILLER_0_283_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13172__B1 _07045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11567__A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15007_ net1221 net1249 game.CPU.applesa.ab.check_walls.above.walls\[35\] vssd1 vssd1
+ vccd1 vccd1 _00225_ sky130_fd_sc_hd__and3_1
X_12219_ _03381_ net421 vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__nor2_1
X_13199_ game.writer.tracker.frame\[400\] game.writer.tracker.frame\[401\] net1023
+ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__mux2_1
XANTENNA__10471__A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_285_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19815_ clknet_leaf_37_clk game.writer.tracker.next_frame\[410\] net1349 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[410\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15981__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16110__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_324_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18707__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__B net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_162_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16958_ net166 _02415_ net91 _02658_ net1496 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[310\]
+ sky130_fd_sc_hd__a32o_1
X_19746_ clknet_leaf_24_clk game.writer.tracker.next_frame\[341\] net1340 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[341\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13475__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_223_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15909_ _01917_ _01918_ _01919_ _01920_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19677_ clknet_leaf_32_clk game.writer.tracker.next_frame\[272\] net1286 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[272\] sky130_fd_sc_hd__dfrtp_1
X_16889_ net145 _02456_ net86 net713 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__o31a_1
XFILLER_0_204_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09430_ net892 net799 game.CPU.applesa.ab.check_walls.above.walls\[114\] net921 vssd1
+ vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__a2bb2o_1
X_18628_ clknet_leaf_8_clk _01045_ _00365_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14424__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16964__A2 _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_301_Right_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09361_ net918 game.CPU.applesa.ab.check_walls.above.walls\[193\] _03485_ net1091
+ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__a22o_1
X_18559_ clknet_leaf_9_clk _00979_ _00296_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11789__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18085__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09292_ net1091 game.CPU.applesa.ab.check_walls.above.walls\[82\] vssd1 vssd1 vccd1
+ vccd1 _03535_ sky130_fd_sc_hd__or2_1
XANTENNA__16177__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload70_A clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10917__Y game.CPU.applesa.ab.absxs.next_head\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_clk_X clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_23 _07032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout131_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__A game.CPU.bad_collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 _02243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_259_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1040_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17141__A2 _02412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10764__A2 _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11961__A1 game.CPU.applesa.ab.check_walls.above.walls\[68\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10652__Y _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12580__B net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16052__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13168__S net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_262_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12910__A0 _06658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1305_A net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11196__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_184_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout765_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19632__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14140__X _08014_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_301_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout932_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14300__B net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09628_ net1139 game.CPU.applesa.ab.absxs.body_y\[18\] vssd1 vssd1 vccd1 vccd1 _03871_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__15115__C game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19782__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16120__A1_N game.CPU.applesa.ab.check_walls.above.walls\[177\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_clk_X clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ net1150 game.CPU.applesa.ab.absxs.body_y\[61\] vssd1 vssd1 vccd1 vccd1 _03802_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_356_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_273_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16508__A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11940__A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12570_ _06442_ _06443_ _06444_ _06446_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__or4b_1
XANTENNA__16168__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12441__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16227__B net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ game.CPU.applesa.ab.check_walls.above.walls\[42\] net768 vssd1 vssd1 vccd1
+ vccd1 _05410_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_137_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11004__X _04894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14240_ game.CPU.applesa.ab.absxs.body_y\[115\] net858 _03323_ net964 vssd1 vssd1
+ vccd1 vccd1 _08114_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11548__A2_N net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11452_ net811 net262 vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10403_ game.CPU.randy.f1.state\[2\] _04341_ _04349_ vssd1 vssd1 vccd1 vccd1 _04552_
+ sky130_fd_sc_hd__and3_1
X_14171_ _08041_ _08042_ _08043_ _08044_ vssd1 vssd1 vccd1 vccd1 _08045_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11383_ net564 _05267_ _05269_ _05271_ _05266_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__o2111a_1
XANTENNA__19650__RESET_B net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17132__A2 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_249_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10755__A2 _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19162__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ game.writer.tracker.frame\[176\] game.writer.tracker.frame\[177\] net1035
+ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__mux2_2
X_10334_ net740 _04490_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__nand2_1
XANTENNA__10562__Y _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_265_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12490__B game.CPU.applesa.twoapples.absxs.next_head\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_284_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13078__S net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13053_ _06923_ _06925_ net687 vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_277_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16891__A1 _02460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17930_ net659 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__inv_2
X_10265_ _04364_ _04365_ _04392_ _04393_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__or4b_1
XANTENNA__11704__A1 game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_226_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1300 net1307 vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__buf_2
XFILLER_0_218_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11704__B2 game.CPU.applesa.ab.check_walls.above.walls\[165\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ _05888_ _05889_ _05890_ _05887_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__a211o_1
Xfanout1311 net1314 vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__buf_2
X_17861_ net2033 _03180_ _03182_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__a21oi_1
Xfanout1322 net1323 vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__buf_2
X_10196_ _04388_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__inv_2
Xfanout1333 net1334 vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__clkbuf_2
Xfanout1344 net1348 vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19600_ clknet_leaf_22_clk game.writer.tracker.next_frame\[195\] net1343 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[195\] sky130_fd_sc_hd__dfrtp_1
Xfanout1355 net1357 vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16643__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16812_ _02499_ net104 net558 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15446__A2 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13457__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17792_ net888 net556 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__nor2_1
Xfanout390 net392 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_2
X_19531_ clknet_leaf_23_clk game.writer.tracker.next_frame\[126\] net1344 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[126\] sky130_fd_sc_hd__dfrtp_1
X_16743_ _02379_ net101 net556 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11834__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13955_ net958 net792 vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__xor2_1
XFILLER_0_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17199__A2 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14413__A2_N net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14210__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19462_ clknet_leaf_40_clk game.writer.tracker.next_frame\[57\] net1358 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[57\] sky130_fd_sc_hd__dfrtp_1
X_12906_ game.writer.tracker.frame\[52\] game.writer.tracker.frame\[53\] net1024 vssd1
+ vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkload7_A clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16674_ net170 _02441_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__nor2_1
X_13886_ net887 game.CPU.applesa.ab.check_walls.above.walls\[96\] net802 net860 _07759_
+ vssd1 vssd1 vccd1 vccd1 _07760_ sky130_fd_sc_hd__a221o_1
XANTENNA__15025__C game.CPU.applesa.ab.check_walls.above.walls\[53\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_271_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18413_ net610 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__inv_2
X_15625_ game.CPU.applesa.ab.check_walls.above.walls\[186\] net465 vssd1 vssd1 vccd1
+ vccd1 _01637_ sky130_fd_sc_hd__xnor2_1
X_12837_ game.writer.tracker.frame\[314\] game.writer.tracker.frame\[315\] net1034
+ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_319_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_295_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19393_ clknet_leaf_55_clk net1397 net1280 vssd1 vssd1 vccd1 vccd1 game.writer.control.detect4.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_319_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12968__A0 _06654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_237_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18344_ net593 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15556_ _08395_ _08926_ _01506_ _01573_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__16159__B1 _01903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12768_ game.writer.tracker.frame\[118\] game.writer.tracker.frame\[119\] net1026
+ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__mux2_1
XANTENNA__12665__B _06507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09320__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14507_ _08377_ _08378_ _08380_ vssd1 vssd1 vccd1 vccd1 _08381_ sky130_fd_sc_hd__or3b_1
XFILLER_0_315_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11719_ net765 _04441_ _04779_ game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1
+ vccd1 vccd1 _05607_ sky130_fd_sc_hd__a31o_1
XANTENNA__15041__B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18275_ net645 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
XANTENNA__13068__S0 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15487_ _01470_ _01511_ _01504_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__o21ai_2
X_12699_ net870 net865 vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__nor2_4
X_17226_ _02542_ net77 _02737_ net1775 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[499\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_13_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19505__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14438_ game.CPU.applesa.ab.absxs.body_x\[88\] net1070 vssd1 vssd1 vccd1 vccd1 _08312_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__14185__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17157_ _02443_ net82 _02718_ game.writer.tracker.frame\[449\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[449\] sky130_fd_sc_hd__a22o_1
XFILLER_0_330_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12681__A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14369_ game.CPU.applesa.ab.absxs.body_y\[117\] net962 vssd1 vssd1 vccd1 vccd1 _08243_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_330_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_326_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16108_ game.CPU.applesa.ab.absxs.body_x\[39\] net461 net440 game.CPU.applesa.ab.absxs.body_y\[38\]
+ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__o22a_1
X_17088_ _02477_ _02692_ _02698_ net1696 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[400\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_283_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_268_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19655__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_248_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16039_ game.CPU.applesa.ab.absxs.body_x\[44\] net271 vssd1 vssd1 vccd1 vccd1 _02051_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_149_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_296_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_271_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16634__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_263_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19729_ clknet_leaf_19_clk game.writer.tracker.next_frame\[324\] net1342 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[324\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13999__A2 game.CPU.applesa.ab.check_walls.above.walls\[74\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_337_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16937__A2 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _03649_ _03650_ _03653_ _03655_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10682__A1 game.CPU.applesa.ab.absxs.body_x\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16328__A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout346_A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11760__A game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09344_ _03581_ _03582_ _03585_ _03586_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__or4_1
XANTENNA__12423__A2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12575__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09230__A game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09275_ net1179 vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout513_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout134_X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1255_A net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19185__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14176__A2 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15886__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17159__A _02237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_X net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_348_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_210_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10737__A2 _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout882_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10823__B _04563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1210_X net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16213__D _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10050_ net1162 _04257_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__nand2_2
XANTENNA__18986__Q game.CPU.applesa.ab.check_walls.above.walls\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11935__A game.CPU.applesa.ab.check_walls.above.walls\[165\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09405__A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_221_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13740_ game.writer.tracker.frame\[245\] game.writer.tracker.frame\[247\] game.writer.tracker.frame\[248\]
+ game.writer.tracker.frame\[246\] net979 net1030 vssd1 vssd1 vccd1 vccd1 _07614_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09899__X _04142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10122__B1 game.CPU.applesa.ab.good_collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ _04834_ _04839_ _04841_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__or3b_1
XANTENNA__16928__A2 _02643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12662__A2 _06531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17050__A1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10673__A1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13671_ net179 _07543_ _07544_ _07542_ vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__o31ai_2
XANTENNA__11870__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ game.CPU.applesa.ab.apple_possible\[4\] net760 game.CPU.applesa.ab.apple_possible\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_195_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15410_ net833 _01430_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__nor2_1
XFILLER_0_183_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15142__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15600__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12622_ _06415_ _06423_ _06485_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__o21a_1
XANTENNA__19528__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16390_ _02252_ net172 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__or2_4
XFILLER_0_38_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10557__Y _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09140__A game.CPU.applesa.ab.check_walls.above.walls\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15341_ game.writer.updater.commands.cmd_num\[2\] _08881_ _08882_ _08877_ vssd1 vssd1
+ vccd1 vccd1 _08883_ sky130_fd_sc_hd__o31a_1
XFILLER_0_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12553_ _03298_ net359 vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11504_ game.CPU.applesa.ab.check_walls.above.walls\[174\] net254 vssd1 vssd1 vccd1
+ vccd1 _05393_ sky130_fd_sc_hd__xnor2_1
X_18060_ net629 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_310_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15272_ _00293_ _08816_ vssd1 vssd1 vccd1 vccd1 _08827_ sky130_fd_sc_hd__nand2_2
XANTENNA__16561__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12484_ _06356_ _06358_ _06359_ _06360_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13375__A0 _06658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_340_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17011_ _02502_ net89 _02674_ net1685 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[347\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18552__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19678__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14223_ game.CPU.applesa.ab.absxs.body_x\[40\] net1073 vssd1 vssd1 vccd1 vccd1 _08097_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__17069__A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_232_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11435_ net777 _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17105__A2 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14154_ net1 _08027_ vssd1 vssd1 vccd1 vccd1 _08028_ sky130_fd_sc_hd__and2_2
X_11366_ game.CPU.applesa.ab.check_walls.above.walls\[34\] net768 vssd1 vssd1 vccd1
+ vccd1 _05255_ sky130_fd_sc_hd__xor2_2
XANTENNA__16864__A1 _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13105_ _06931_ _06932_ net682 vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_238_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10317_ game.CPU.randy.f1.a1.count\[14\] _04495_ vssd1 vssd1 vccd1 vccd1 _04499_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_237_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11297_ _04877_ _04879_ _04880_ _04881_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__or4_1
X_18962_ net1200 _00265_ _00633_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_14085_ _03374_ net807 net805 net854 _07955_ vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__a221o_1
XFILLER_0_265_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13036_ net681 _06891_ _06909_ net506 vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__o211a_1
XFILLER_0_253_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10248_ net779 net771 vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__and2_4
X_17913_ net662 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__inv_2
XFILLER_0_237_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18893_ clknet_leaf_2_clk _01265_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_266_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1130 net1133 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__buf_4
Xfanout1141 net1143 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__buf_2
X_17844_ _03169_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_321_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10179_ _04366_ _04371_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__xnor2_1
Xfanout1152 game.CPU.applesa.ab.snake_head_y\[1\] vssd1 vssd1 vccd1 vccd1 net1152
+ sky130_fd_sc_hd__buf_4
XFILLER_0_266_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1163 net1165 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_4
Xfanout1174 game.CPU.applesa.ab.XMAX\[2\] vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__buf_2
XFILLER_0_206_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1185 net1186 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__buf_2
XANTENNA__09315__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19058__CLK net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17775_ game.CPU.applesa.twoapples.count\[0\] net1163 vssd1 vssd1 vccd1 vccd1 _03126_
+ sky130_fd_sc_hd__nor2_1
Xfanout1196 net1198 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__clkbuf_2
X_14987_ net1225 net1252 game.CPU.applesa.ab.check_walls.above.walls\[15\] vssd1 vssd1
+ vccd1 vccd1 _00203_ sky130_fd_sc_hd__and3_1
XFILLER_0_282_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16726_ _02359_ _02561_ net735 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__o21a_1
X_19514_ clknet_leaf_28_clk game.writer.tracker.next_frame\[109\] net1283 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[109\] sky130_fd_sc_hd__dfrtp_1
X_13938_ _07807_ _07808_ _07811_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__or3_1
XANTENNA__13850__A1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12653__A2 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16919__A2 _02643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13850__B2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17041__A1 _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17041__B2 game.writer.tracker.frame\[368\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19445_ clknet_leaf_47_clk game.writer.tracker.next_frame\[40\] net1298 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[40\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_347_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16657_ net190 net128 _02418_ _02547_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[120\]
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_85_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12676__A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13869_ game.CPU.applesa.ab.XMAX\[0\] net886 net1060 _03370_ vssd1 vssd1 vccd1 vccd1
+ _07743_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_201_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15608_ game.CPU.applesa.ab.absxs.body_y\[34\] net333 vssd1 vssd1 vccd1 vccd1 _01620_
+ sky130_fd_sc_hd__or2_1
X_19376_ clknet_leaf_9_clk _01382_ _00957_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.snake_head_y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_16588_ net171 net151 _02348_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09806__B1 game.CPU.applesa.ab.check_walls.above.walls\[106\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_335_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09050__A game.CPU.applesa.ab.absxs.body_y\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18327_ net599 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15539_ _01492_ _01512_ _01538_ _01560_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_157_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_332_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19572__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_301_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09060_ game.CPU.applesa.ab.absxs.body_y\[46\] vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__inv_2
XANTENNA__14158__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18258_ net622 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_170_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13366__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17209_ net146 _02369_ net75 _02733_ net1479 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[486\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12169__B2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18189_ net609 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__inv_2
XANTENNA__10483__X _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10924__A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold602 game.writer.tracker.frame\[408\] vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11916__A1 game.CPU.applesa.ab.check_walls.above.walls\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10719__A2 _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold613 game.CPU.applesa.ab.count_luck\[1\] vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold624 game.CPU.clock1.counter\[13\] vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11739__B net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold635 game.CPU.walls.rand_wall.inputa vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload33_A clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold646 game.CPU.apple_location\[3\] vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 game.writer.tracker.frame\[337\] vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16855__B2 game.writer.tracker.frame\[241\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold668 game.CPU.applesa.ab.absxs.body_y\[25\] vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ net1261 game.CPU.bodymain1.Direction\[0\] vssd1 vssd1 vccd1 vccd1 _04192_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__16611__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14330__A2 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09893_ _03748_ _04085_ _04134_ _04135_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_168_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16330__B _02322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_271_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout296_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_181_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14131__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1003_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17280__A1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09225__A game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__B net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout463_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15514__X net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12644__A2 _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16329__Y _02322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17032__A1 _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10655__A1 game.CPU.applesa.ab.absxs.body_x\[35\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_X net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10655__B2 game.CPU.applesa.ab.absxs.body_x\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout728_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_342_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_270_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_260_Left_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09327_ net910 game.CPU.applesa.ab.absxs.body_x\[80\] _03330_ net1144 _03569_ vssd1
+ vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12947__A3 _06813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18273__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1160_X net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19820__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ game.CPU.randy.counter1.count\[7\] vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_322_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09189_ game.CPU.applesa.ab.check_walls.above.walls\[108\] vssd1 vssd1 vccd1 vccd1
+ _03438_ sky130_fd_sc_hd__inv_2
XFILLER_0_279_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_177_Right_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14306__A game.CPU.applesa.ab.absxs.body_x\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11907__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17099__A1 _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11220_ _03245_ net413 vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nand2_1
XANTENNA__11907__B2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_294_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11649__B game.CPU.applesa.ab.apple_possible\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19970__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14025__B game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_268_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10040__C1 game.CPU.applesa.ab.YMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11151_ game.CPU.applesa.ab.absxs.body_y\[99\] net400 net414 game.CPU.applesa.ab.absxs.body_x\[97\]
+ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__15649__A2 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_281_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10102_ net846 _04305_ _04309_ net1271 vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__a22o_1
XANTENNA__14321__A2 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11082_ _04970_ _04971_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__nor2_1
XANTENNA__13755__S1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19605__Q game.writer.tracker.frame\[200\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19200__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14910_ net1170 _08428_ _08430_ net1174 _08686_ vssd1 vssd1 vccd1 vccd1 _08687_ sky130_fd_sc_hd__o221a_1
X_10033_ _04236_ _04240_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__nand2_1
XANTENNA__11665__A game.CPU.applesa.ab.check_walls.above.walls\[121\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15137__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15890_ _01898_ _01899_ _01900_ _01901_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_145_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17271__A1 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09135__A game.CPU.applesa.ab.check_walls.above.walls\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14841_ game.CPU.randy.f1.c1.count\[3\] game.CPU.randy.f1.c1.count\[4\] _08632_ game.CPU.randy.f1.c1.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _08640_ sky130_fd_sc_hd__a31o_1
XANTENNA__14085__A1 _03374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_230_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18448__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14085__B2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17560_ _02879_ _02918_ _02939_ _02985_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__or4_1
XANTENNA__12096__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14772_ game.CPU.randy.counter1.count\[12\] game.CPU.randy.counter1.count\[11\] net265
+ vssd1 vssd1 vccd1 vccd1 _08593_ sky130_fd_sc_hd__a21o_1
XANTENNA__19350__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ net784 net554 vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__or2_1
X_16511_ net221 _02453_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__nor2_8
XTAP_TAPCELL_ROW_205_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13723_ game.writer.tracker.frame\[194\] net843 net837 game.writer.tracker.frame\[193\]
+ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__o22a_1
XFILLER_0_357_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10935_ _03291_ net412 vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__nand2_1
X_17491_ net846 _02778_ net428 _02919_ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__a31o_1
XANTENNA__18918__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19230_ clknet_leaf_57_clk net1424 _00868_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.normal1.number\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_292_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16442_ net196 _02399_ _02402_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__a21o_4
XFILLER_0_183_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_357_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_317_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13045__C1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13654_ game.writer.tracker.frame\[5\] game.writer.tracker.frame\[7\] game.writer.tracker.frame\[8\]
+ game.writer.tracker.frame\[6\] net969 net1005 vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14388__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_clk_X clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10866_ game.CPU.randy.counter1.count\[6\] _03508_ game.CPU.randy.counter1.count\[5\]
+ _03510_ _04744_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_234_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ game.CPU.applesa.ab.absxs.body_y\[62\] net521 net365 net1270 _06481_ vssd1
+ vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__a221o_1
XFILLER_0_183_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19161_ clknet_leaf_70_clk _00290_ _00832_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.input2
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16373_ net1979 net734 _02352_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[31\]
+ sky130_fd_sc_hd__and3_1
X_13585_ game.writer.tracker.frame\[338\] net843 net675 game.writer.tracker.frame\[340\]
+ _07458_ vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__o221a_1
XANTENNA__17326__A2 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10797_ game.CPU.applesa.ab.absxs.body_y\[40\] _04690_ _04728_ game.CPU.applesa.ab.absxs.body_y\[36\]
+ vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__a22o_1
X_18112_ net583 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__inv_2
XANTENNA__10949__A2 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10447__C net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15324_ _08868_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19092_ net1178 _00129_ _00763_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[137\]
+ sky130_fd_sc_hd__dfrtp_4
X_12536_ game.CPU.applesa.ab.absxs.body_y\[42\] net519 vssd1 vssd1 vccd1 vccd1 _06413_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_23_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13348__A0 _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18043_ net659 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_312_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15255_ game.CPU.kyle.L1.nextState\[3\] _08809_ net264 net1877 vssd1 vssd1 vccd1
+ vccd1 _01264_ sky130_fd_sc_hd__a22o_2
X_12467_ game.CPU.applesa.ab.absxs.body_x\[14\] net372 vssd1 vssd1 vccd1 vccd1 _06344_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10744__A game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14206_ game.CPU.applesa.ab.absxs.body_x\[67\] net875 net865 game.CPU.applesa.ab.absxs.body_y\[65\]
+ _08077_ vssd1 vssd1 vccd1 vccd1 _08080_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_285_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11418_ net743 _05302_ _05305_ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__a211o_1
XANTENNA__11559__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15186_ _08755_ _08757_ vssd1 vssd1 vccd1 vccd1 _08761_ sky130_fd_sc_hd__and2b_1
X_12398_ game.CPU.applesa.ab.absxs.body_y\[92\] net359 vssd1 vssd1 vccd1 vccd1 _06275_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10463__B _04594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11374__A2 _05207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14137_ net1070 _03401_ game.CPU.applesa.ab.check_walls.above.walls\[41\] net882
+ vssd1 vssd1 vccd1 vccd1 _08011_ sky130_fd_sc_hd__a22o_1
X_11349_ net742 _05235_ _05236_ net563 vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__a2bb2o_1
X_19994_ clknet_leaf_45_clk _01418_ net1299 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_245_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14312__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14068_ net945 net831 vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__xnor2_1
X_18945_ net1175 _00084_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number_out\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12323__A1 _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13019_ _06877_ _06878_ net485 vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18876_ clknet_leaf_5_clk game.CPU.randy.f1.c1.innerCount\[6\] _00571_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17262__A1 _02275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10885__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09045__A game.CPU.applesa.ab.absxs.body_y\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17827_ game.writer.updater.commands.count\[4\] game.writer.updater.commands.count\[3\]
+ _03153_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__and3_1
XFILLER_0_240_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14076__A1 game.CPU.applesa.ab.YMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_233_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14886__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15812__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13823__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17758_ net1902 _03113_ _03114_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_334_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10637__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16709_ _02238_ net140 net559 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a21oi_2
XANTENNA__18598__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17689_ game.CPU.walls.rand_wall.count_luck\[4\] _03068_ net1976 vssd1 vssd1 vccd1
+ vccd1 _03072_ sky130_fd_sc_hd__a21oi_1
XANTENNA__19843__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_279_Right_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15603__A2_N net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19428_ clknet_leaf_41_clk game.writer.tracker.next_frame\[23\] net1331 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[23\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13036__C1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10638__B _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19359_ clknet_leaf_68_clk _01365_ _00940_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_29_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17317__A2 _02416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13682__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_350_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09112_ net1274 vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_98_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19993__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_304_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16325__B _02318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09043_ game.CPU.applesa.ab.absxs.body_x\[8\] vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14000__A1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout211_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10654__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14000__B2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_A _05606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold410 game.writer.tracker.frame\[538\] vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_345_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold421 game.writer.tracker.frame\[520\] vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 game.writer.tracker.frame\[197\] vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 game.writer.tracker.frame\[459\] vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19223__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold454 game.writer.tracker.frame\[319\] vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold465 game.writer.tracker.frame\[575\] vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 game.writer.tracker.frame\[361\] vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 game.writer.tracker.frame\[481\] vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1218_A game.CPU.walls.rand_wall.start_enable vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold498 game.writer.tracker.frame\[54\] vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 _03201_ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_4
XFILLER_0_256_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14303__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09945_ _04180_ _04181_ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__and2_1
Xfanout912 net913 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout580_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout923 _03193_ vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_229_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout934 net935 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16060__B net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout678_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net946 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__buf_2
XANTENNA_fanout299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13511__B1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_256_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11485__A game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net957 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_216_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout967 net972 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__buf_4
X_09876_ _04050_ _04053_ _03704_ _04016_ _04042_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__o2111a_1
Xfanout978 net979 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__buf_4
XANTENNA__19373__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16995__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout989 net994 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__buf_2
XANTENNA__17253__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16056__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09730__A2 game.CPU.applesa.ab.absxs.body_x\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout845_A _06574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18268__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12617__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_356_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17005__A1 _02491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12587__Y _06464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11932__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_246_Right_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17900__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10720_ game.CPU.applesa.ab.absxs.body_y\[46\] _04640_ _04641_ game.CPU.applesa.ab.absxs.body_y\[42\]
+ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__a22o_1
XFILLER_0_339_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15123__C net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13578__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _04694_ game.CPU.applesa.ab.absxs.body_x\[40\] _04690_ vssd1 vssd1 vccd1
+ vccd1 _01111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16516__A _02267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13673__S0 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13370_ _06683_ _06685_ net693 vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__mux2_1
X_10582_ game.CPU.applesa.ab.absxs.body_x\[115\] _04663_ _04664_ game.CPU.applesa.ab.absxs.body_x\[111\]
+ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_307_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_298_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10800__A1 game.CPU.applesa.ab.absxs.body_y\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12321_ _06129_ _06131_ _06132_ _06157_ _06091_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__o311a_1
XFILLER_0_145_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16531__A3 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15040_ net1219 net1248 game.CPU.applesa.ab.check_walls.above.walls\[68\] vssd1 vssd1
+ vccd1 vccd1 _00261_ sky130_fd_sc_hd__and3_1
XFILLER_0_310_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11379__B net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ net803 net419 vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_279_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16819__A1 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11203_ game.CPU.applesa.ab.absxs.body_y\[92\] net533 vssd1 vssd1 vccd1 vccd1 _05093_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__13875__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12183_ _05935_ _06068_ _05937_ _05936_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__or4bb_1
XANTENNA_clkbuf_leaf_61_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16251__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19716__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16295__A2 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ game.CPU.applesa.ab.absxs.body_y\[69\] net542 vssd1 vssd1 vccd1 vccd1 _05024_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_275_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16991_ _02472_ net88 _02668_ net1736 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[333\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17066__B _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_247_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18730_ clknet_leaf_13_clk _01147_ _00467_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[112\]
+ sky130_fd_sc_hd__dfrtp_4
X_11065_ _03350_ net405 vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__xnor2_1
X_15942_ _03404_ net332 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__nor2_1
XANTENNA__09136__Y _03385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17244__A1 _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ net1163 game.CPU.applesa.out_random_2\[3\] vssd1 vssd1 vccd1 vccd1 _04224_
+ sky130_fd_sc_hd__nand2_1
X_18661_ clknet_leaf_60_clk _01078_ _00398_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[79\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_222_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15873_ game.CPU.applesa.ab.absxs.body_y\[24\] net451 vssd1 vssd1 vccd1 vccd1 _01885_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_215_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18740__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15255__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13814__S net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19866__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14824_ net139 _08628_ _08629_ vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__and3_1
X_17612_ net1860 _03021_ net429 vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_240_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18592_ clknet_leaf_50_clk _01012_ _00329_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[65\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_24_Left_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_230_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17543_ _03219_ game.CPU.speed1.Qa\[0\] net426 _02936_ _02958_ vssd1 vssd1 vccd1
+ vccd1 _02970_ sky130_fd_sc_hd__a311o_1
X_14755_ game.CPU.randy.counter1.count1\[17\] _08575_ vssd1 vssd1 vccd1 vccd1 _08578_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09485__A1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19070__Q game.CPU.applesa.ab.check_walls.above.walls\[115\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ _05617_ _05636_ _05711_ _05854_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.collision_rightn
+ sky130_fd_sc_hd__or4_1
XANTENNA__17547__A2 game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09485__B2 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ net209 _07579_ vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13018__C1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10918_ game.CPU.applesa.ab.logic_enable net846 net1272 vssd1 vssd1 vccd1 vccd1 _04813_
+ sky130_fd_sc_hd__a21oi_1
X_17474_ _02889_ _02897_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_213_Right_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15033__C game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14686_ _08503_ _08523_ _08524_ vssd1 vssd1 vccd1 vccd1 _08525_ sky130_fd_sc_hd__o21ba_1
X_11898_ net573 _05409_ _05410_ net751 vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__a22o_1
XFILLER_0_345_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16425_ net135 net115 _02390_ _02388_ net1481 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[45\]
+ sky130_fd_sc_hd__a32o_1
X_19213_ net1169 _00025_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_possible\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_13637_ game.writer.tracker.frame\[17\] game.writer.tracker.frame\[19\] game.writer.tracker.frame\[20\]
+ game.writer.tracker.frame\[18\] net977 net1024 vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10849_ _03506_ game.CPU.randy.counter1.count1\[7\] _03505_ game.CPU.randy.counter1.count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__16426__A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19144_ net1187 _00186_ _00815_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[189\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16356_ net197 _02340_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__nor2_4
XANTENNA_clkbuf_leaf_14_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16507__B1 _02450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13568_ game.writer.tracker.frame\[329\] game.writer.tracker.frame\[331\] game.writer.tracker.frame\[332\]
+ game.writer.tracker.frame\[330\] net968 net998 vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__mux4_1
XANTENNA__16145__B net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15307_ game.CPU.applesa.twomode.number\[3\] _08849_ vssd1 vssd1 vccd1 vccd1 _08854_
+ sky130_fd_sc_hd__or2_1
X_12519_ game.CPU.applesa.ab.absxs.body_x\[69\] net379 vssd1 vssd1 vccd1 vccd1 _06396_
+ sky130_fd_sc_hd__nor2_1
X_19075_ net1179 _00111_ _00746_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[120\]
+ sky130_fd_sc_hd__dfrtp_4
X_16287_ net244 _02227_ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13499_ _07067_ _07069_ _07073_ _07068_ net705 net497 vssd1 vssd1 vccd1 vccd1 _07373_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__17180__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_251_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_301_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18026_ net662 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__inv_2
X_15238_ net577 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__inv_2
XFILLER_0_313_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15984__B net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13741__A0 game.writer.tracker.frame\[241\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15169_ net1227 net1254 game.CPU.walls.rand_wall.y_final\[1\] vssd1 vssd1 vccd1 vccd1
+ _00243_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_93_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout208 net218 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_4
Xfanout219 net223 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_4
X_19977_ clknet_leaf_39_clk game.writer.tracker.next_frame\[572\] net1330 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[572\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14297__A1 game.CPU.applesa.ab.absxs.body_x\[55\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_266_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_238_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09730_ net921 game.CPU.applesa.ab.absxs.body_x\[34\] _03347_ net1155 _03972_ vssd1
+ vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__a221o_1
X_18928_ clknet_leaf_6_clk net3 _00612_ vssd1 vssd1 vccd1 vccd1 game.CPU.right_button.sync1.Q
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_348_Right_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_165_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_340_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09661_ net1084 _03243_ game.CPU.applesa.ab.absxs.body_x\[38\] net922 vssd1 vssd1
+ vccd1 vccd1 _03904_ sky130_fd_sc_hd__a22o_1
X_18859_ clknet_leaf_1_clk _01250_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__19934__RESET_B net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18088__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15505__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09592_ _03831_ _03832_ _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__or3b_1
XFILLER_0_221_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout259_A _05195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_323_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12480__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_336_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1070_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16336__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13655__S0 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_351_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16761__A3 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12583__B net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1335_A net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19739__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18613__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09026_ game.CPU.applesa.ab.absxs.body_x\[34\] vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__inv_2
XANTENNA__15894__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13732__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold240 game.writer.tracker.frame\[358\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 game.writer.tracker.frame\[439\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14143__X _08017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1123_X net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09400__A1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold262 game.writer.tracker.frame\[562\] vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09400__B2 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold273 game.writer.tracker.frame\[426\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_265_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_348_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold284 game.writer.tracker.frame\[274\] vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 game.writer.tracker.frame\[356\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_207_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_291_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_244_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout962_A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_272_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout720 net721 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__buf_2
XANTENNA__18763__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout731 net738 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__clkbuf_2
XANTENNA__19889__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_187_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout742 _04451_ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__buf_4
X_09928_ net1100 net1262 _04158_ _04167_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_315_Right_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout764 game.CPU.applesa.ab.apple_possible\[3\] vssd1 vssd1 vccd1 vccd1 net764
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout74_A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17226__A1 _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14121__A2_N net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout775 net776 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_304_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout786 game.CPU.applesa.ab.check_walls.above.walls\[167\] vssd1 vssd1 vccd1 vccd1
+ net786 sky130_fd_sc_hd__clkbuf_4
X_20048_ game.CPU.kyle.L1.lcd_rs vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XANTENNA__18994__Q game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_272_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09859_ net1086 game.CPU.applesa.ab.absxs.body_x\[47\] vssd1 vssd1 vccd1 vccd1 _04102_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_6_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout797 game.CPU.applesa.ab.check_walls.above.walls\[118\] vssd1 vssd1 vccd1 vccd1
+ net797 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12870_ game.writer.tracker.frame\[40\] game.writer.tracker.frame\[41\] net992 vssd1
+ vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_358_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11662__B net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11821_ _05701_ _05702_ _05708_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__or3_1
XFILLER_0_200_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15134__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_202_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_276_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _08407_ _08411_ _08412_ net556 vssd1 vssd1 vccd1 vccd1 game.writer.control.next\[1\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_212_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11752_ net569 _05388_ _05383_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_218_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ game.CPU.applesa.ab.absxs.body_y\[71\] _04625_ _04626_ game.CPU.applesa.ab.absxs.body_y\[67\]
+ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__a22o_1
XANTENNA__19269__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14471_ _08337_ _08338_ _08340_ _08344_ vssd1 vssd1 vccd1 vccd1 _08345_ sky130_fd_sc_hd__or4_2
XFILLER_0_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11683_ game.CPU.applesa.ab.check_walls.above.walls\[56\] net778 vssd1 vssd1 vccd1
+ vccd1 _05572_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_354_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13222__X _07096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16752__A3 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16210_ _01605_ _02219_ _02221_ _01976_ _01597_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__o2111a_4
X_13422_ net696 _06995_ _07295_ net504 vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__o211a_1
XANTENNA__15150__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17190_ net149 _02497_ net77 _02728_ net1674 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[472\]
+ sky130_fd_sc_hd__a32o_1
X_10634_ _03271_ net561 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11577__A2 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16141_ game.CPU.applesa.ab.absxs.body_x\[78\] net347 vssd1 vssd1 vccd1 vccd1 _02153_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_342_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13353_ _06640_ _06650_ _06652_ _06651_ net510 net703 vssd1 vssd1 vccd1 vccd1 _07227_
+ sky130_fd_sc_hd__mux4_1
X_10565_ game.CPU.applesa.ab.absxs.body_x\[14\] _04653_ _04654_ game.CPU.applesa.ab.absxs.body_x\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12304_ _03405_ net421 vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__nor2_1
XANTENNA__14515__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16072_ game.CPU.applesa.ab.absxs.body_y\[85\] net444 vssd1 vssd1 vccd1 vccd1 _02084_
+ sky130_fd_sc_hd__xnor2_1
X_13284_ _07156_ _07157_ net487 vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17348__Y _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10496_ _04177_ _04614_ _04618_ _04578_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__a31o_1
XFILLER_0_295_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13723__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_258_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19900_ clknet_leaf_15_clk game.writer.tracker.next_frame\[495\] net1288 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[495\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14153__D_N _08026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15023_ net1222 net1250 game.CPU.applesa.ab.check_walls.above.walls\[51\] vssd1 vssd1
+ vccd1 vccd1 _00242_ sky130_fd_sc_hd__and3_1
XFILLER_0_310_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12235_ game.CPU.applesa.ab.check_walls.above.walls\[71\] net424 vssd1 vssd1 vccd1
+ vccd1 _06121_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_287_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10537__B1 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19831_ clknet_leaf_33_clk game.writer.tracker.next_frame\[426\] net1325 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[426\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_229_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12166_ game.CPU.applesa.ab.check_walls.above.walls\[156\] net552 vssd1 vssd1 vccd1
+ vccd1 _06053_ sky130_fd_sc_hd__or2_1
XANTENNA__14213__B net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13892__X _07766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_242_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ game.CPU.applesa.ab.absxs.body_y\[19\] net397 vssd1 vssd1 vccd1 vccd1 _05007_
+ sky130_fd_sc_hd__xnor2_1
X_19762_ clknet_leaf_30_clk game.writer.tracker.next_frame\[357\] net1292 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[357\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17805__A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16974_ _02450_ net90 _02662_ net1784 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[322\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13487__C1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ net803 net290 net296 net802 vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__17217__A1 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18713_ clknet_leaf_52_clk _01130_ _00450_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[75\]
+ sky130_fd_sc_hd__dfrtp_4
X_15925_ _01925_ _01926_ _01932_ _01933_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__or4_1
X_11048_ _03330_ net405 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__xnor2_2
X_19693_ clknet_leaf_26_clk game.writer.tracker.next_frame\[288\] net1313 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[288\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_274_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput8 nrst vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_1
X_15856_ game.CPU.applesa.ab.absxs.body_x\[99\] net458 net445 game.CPU.applesa.ab.absxs.body_y\[97\]
+ _01861_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a221o_1
X_18644_ clknet_leaf_53_clk _01061_ _00381_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[46\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_349_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_318_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14807_ net1662 _08616_ _08618_ vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11572__B net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09458__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18575_ clknet_leaf_61_clk _00995_ _00312_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[32\]
+ sky130_fd_sc_hd__dfrtp_4
X_15787_ game.CPU.applesa.ab.absxs.body_x\[75\] net460 vssd1 vssd1 vccd1 vccd1 _01799_
+ sky130_fd_sc_hd__xnor2_1
X_12999_ game.writer.tracker.frame\[530\] game.writer.tracker.frame\[531\] net1007
+ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__mux2_1
XANTENNA__09458__B2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11349__A1_N net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17526_ game.CPU.kyle.L1.nextState\[0\] _04484_ _02835_ _04482_ vssd1 vssd1 vccd1
+ vccd1 _02954_ sky130_fd_sc_hd__o211a_1
X_14738_ _08565_ _08566_ net55 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__and3b_1
XANTENNA__15979__B net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10188__B net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17457_ _04638_ _02784_ _02789_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14669_ game.CPU.randy.counter1.count1\[7\] _08498_ vssd1 vssd1 vccd1 vccd1 _08508_
+ sky130_fd_sc_hd__and2_1
XANTENNA__13637__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12684__A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_313_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16408_ net163 _02377_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__and2_4
XFILLER_0_333_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18636__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13411__C1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17388_ _02816_ _02817_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_41_Left_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16339_ net134 _02259_ _02328_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__or3_1
X_19127_ net1183 _00168_ _00798_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[172\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09630__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09630__B2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_301_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19058_ net1194 _00092_ _00729_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_298_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14506__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_329_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18786__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18009_ net643 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__inv_2
XFILLER_0_301_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10528__B1 _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__A game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_168_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16322__C _06607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09713_ net1109 game.CPU.applesa.ab.absxs.body_x\[20\] vssd1 vssd1 vccd1 vccd1 _03956_
+ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout376_A _06209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_260_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09644_ net1089 _03459_ _03460_ net1082 vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_3_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09449__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09575_ net1098 _03402_ _03403_ net1146 vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a22o_1
XANTENNA__19411__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09449__B2 net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_353_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17450__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16719__B1 _02574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15889__B net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13650__C1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout710_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_336_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout808_A game.CPU.applesa.ab.check_walls.above.walls\[87\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_X net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19561__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_324_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1240_X net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18281__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11964__C1 _05830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_213_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18989__Q game.CPU.applesa.ab.check_walls.above.walls\[34\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10350_ game.CPU.walls.rand_wall.counter2\[4\] game.CPU.walls.rand_wall.counter2\[3\]
+ game.CPU.walls.rand_wall.counter2\[1\] vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_189_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16513__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13629__S net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ game.CPU.applesa.ab.absxs.body_x\[110\] vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__inv_2
X_10281_ net851 game.CPU.applesa.ab.good_spot_next vssd1 vssd1 vccd1 vccd1 _04473_
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_3_0_clk_X clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _05904_ _05905_ _05906_ _05903_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__a211o_1
XANTENNA__09408__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__B net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout965_X net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout77_X net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 _04786_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_4
Xfanout561 net562 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_2
Xfanout572 net575 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_2
Xfanout583 net585 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_4
X_13971_ net1054 game.CPU.applesa.ab.check_walls.above.walls\[82\] vssd1 vssd1 vccd1
+ vccd1 _07845_ sky130_fd_sc_hd__xnor2_1
Xfanout594 net595 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_4
XANTENNA__13364__S net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15710_ _03290_ net348 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11673__A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ _06696_ _06698_ net678 vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__mux2_1
XANTENNA__15145__A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16690_ _02466_ net62 _02563_ net1962 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[137\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_224_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12488__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16422__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09143__A game.CPU.applesa.ab.check_walls.above.walls\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15641_ _03265_ net346 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11392__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ game.writer.tracker.frame\[270\] game.writer.tracker.frame\[271\] net996
+ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_347_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14984__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_319_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15630__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18360_ net597 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__inv_2
X_11804_ game.CPU.applesa.ab.check_walls.above.walls\[61\] net308 vssd1 vssd1 vccd1
+ vccd1 _05692_ sky130_fd_sc_hd__or2_1
XANTENNA__12444__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15572_ net1431 net1429 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__xnor2_1
XANTENNA__18659__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12784_ game.writer.tracker.frame\[352\] game.writer.tracker.frame\[353\] net1013
+ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__mux2_1
XANTENNA__19904__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17311_ net130 _02535_ net1647 net724 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[562\]
+ sky130_fd_sc_hd__o211a_1
X_14523_ _07400_ _07742_ _08396_ _07164_ vssd1 vssd1 vccd1 vccd1 _08397_ sky130_fd_sc_hd__o31ai_1
XANTENNA__11798__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11735_ net801 net301 _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__o21ba_1
X_18291_ net623 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
XANTENNA__13619__S0 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20009__1378 vssd1 vssd1 vccd1 vccd1 net1378 _20009__1378/LO sky130_fd_sc_hd__conb_1
XANTENNA__16186__B2 game.CPU.applesa.ab.check_walls.above.walls\[106\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17242_ _02552_ net79 _02741_ net1781 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[511\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_327_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14454_ _03319_ net964 net946 _03318_ vssd1 vssd1 vccd1 vccd1 _08328_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11666_ net774 _05554_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_289_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ net680 _06867_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17173_ _02470_ net73 _02724_ net1828 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[459\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13944__B1 game.CPU.applesa.ab.check_walls.above.walls\[70\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10617_ game.CPU.applesa.ab.absxs.body_x\[72\] _04675_ _04676_ game.CPU.applesa.ab.absxs.body_x\[68\]
+ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17135__B1 _02713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09612__A1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14385_ game.CPU.applesa.ab.absxs.body_y\[4\] net869 _03225_ net1063 vssd1 vssd1
+ vccd1 vccd1 _08259_ sky130_fd_sc_hd__a2bb2o_1
X_11597_ _05483_ _05484_ _05485_ _05482_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__and4b_1
XANTENNA__09612__B2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16124_ _03465_ net350 net465 game.CPU.applesa.ab.check_walls.above.walls\[162\]
+ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__a22o_1
X_13336_ _06611_ _06621_ _06625_ _06624_ net501 net693 vssd1 vssd1 vccd1 vccd1 _07210_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10548_ net850 _04644_ _04646_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__or3b_2
XFILLER_0_134_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_269_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15697__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11848__A game.CPU.applesa.ab.check_walls.above.walls\[53\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16055_ _02062_ _02064_ _02065_ _02066_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__or4_1
XFILLER_0_295_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13267_ _07139_ _07140_ net479 vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__mux2_1
X_10479_ _04358_ _04578_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__nor2_8
XANTENNA__13172__A1 _07000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15006_ net1220 net1248 game.CPU.applesa.ab.check_walls.above.walls\[34\] vssd1 vssd1
+ vccd1 vccd1 _00224_ sky130_fd_sc_hd__and3_1
XANTENNA__13172__B2 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09318__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ game.CPU.applesa.ab.check_walls.above.walls\[6\] net420 vssd1 vssd1 vccd1
+ vccd1 _06104_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11567__B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13198_ net242 _07059_ _07071_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__or3_1
XANTENNA__11722__A2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19814_ clknet_leaf_37_clk game.writer.tracker.next_frame\[409\] net1349 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[409\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16110__A1 game.CPU.applesa.ab.check_walls.above.walls\[11\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ net793 net551 vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__nand2_1
XFILLER_0_208_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_324_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14121__B1 game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16661__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19745_ clknet_leaf_24_clk game.writer.tracker.next_frame\[340\] net1340 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[340\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_236_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16957_ _02412_ net94 _02658_ net1617 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[309\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19434__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13274__S net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11583__A _05423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15908_ game.CPU.applesa.ab.absxs.body_x\[58\] net467 vssd1 vssd1 vccd1 vccd1 _01920_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__11486__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19676_ clknet_leaf_32_clk game.writer.tracker.next_frame\[271\] net1286 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[271\] sky130_fd_sc_hd__dfrtp_1
X_16888_ _02241_ net120 vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__nand2_4
XANTENNA__12398__B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09053__A game.CPU.applesa.ab.absxs.body_y\[76\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18627_ clknet_leaf_16_clk _01044_ _00364_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_0_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10199__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15839_ game.CPU.applesa.ab.check_walls.above.walls\[19\] net462 vssd1 vssd1 vccd1
+ vccd1 _01851_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12966__X _06840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14894__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_304_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13858__S0 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09360_ net1147 game.CPU.applesa.ab.check_walls.above.walls\[197\] vssd1 vssd1 vccd1
+ vccd1 _03603_ sky130_fd_sc_hd__xor2_1
XANTENNA__19584__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18558_ clknet_leaf_1_clk _00014_ _00295_ vssd1 vssd1 vccd1 vccd1 game.CPU.speed1.Qa\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17509_ _02853_ _02920_ _02922_ _02935_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__or4_1
X_09291_ net1156 net810 vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__or2_1
X_18489_ net583 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__inv_2
XANTENNA__16177__B2 game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_13 _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_24 _07032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_35 _07620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_46 _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload63_A clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16614__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout124_A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_259_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_259_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17141__A3 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16333__B net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11961__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1033_A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13699__C1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14360__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09228__A game.CPU.applesa.ab.check_walls.above.walls\[179\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_262_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1200_A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_184_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout660_A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_301_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_345_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11477__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13871__C1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19927__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09627_ net1130 game.CPU.applesa.ab.absxs.body_y\[19\] vssd1 vssd1 vccd1 vccd1 _03870_
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1190_X net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout925_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12101__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18276__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09558_ _03797_ _03798_ _03799_ _03800_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__or4b_1
XFILLER_0_210_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_273_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16508__B _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18951__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ net1106 game.CPU.applesa.ab.check_walls.above.walls\[184\] vssd1 vssd1 vccd1
+ vccd1 _03732_ sky130_fd_sc_hd__xor2_1
XFILLER_0_92_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ game.CPU.applesa.ab.check_walls.above.walls\[43\] net763 vssd1 vssd1 vccd1
+ vccd1 _05409_ sky130_fd_sc_hd__xnor2_2
XANTENNA__15131__C net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11451_ _05335_ _05337_ _05339_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__and3_1
XANTENNA__17117__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10402_ game.CPU.randy.f1.state\[4\] _04550_ _04551_ vssd1 vssd1 vccd1 vccd1 _01244_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_351_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14170_ game.CPU.applesa.ab.absxs.body_y\[105\] net964 vssd1 vssd1 vccd1 vccd1 _08044_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11401__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11382_ net564 _05267_ _05265_ net743 vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__20046__A game.CPU.randy.counter1.out vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17132__A3 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13359__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13121_ game.writer.tracker.frame\[172\] game.writer.tracker.frame\[173\] net990
+ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10333_ net740 _04489_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__nand2_1
XFILLER_0_249_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14044__A net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13052_ game.writer.tracker.frame\[254\] game.writer.tracker.frame\[255\] net1032
+ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_284_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11387__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10264_ _04455_ _04456_ net1173 _03493_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11165__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19457__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16530__Y _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_226_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12003_ _05584_ _05586_ _05587_ _05589_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__or4_1
XANTENNA__11704__A2 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11955__X _05843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1301 net1302 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17355__A _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13883__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1312 net1313 vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__clkbuf_4
X_17860_ game.writer.updater.commands.count\[13\] _03180_ _03175_ vssd1 vssd1 vccd1
+ vccd1 _03182_ sky130_fd_sc_hd__o21ai_1
X_10195_ _04382_ _04387_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__and2_1
Xfanout1323 net1360 vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__clkbuf_2
Xfanout1334 net1360 vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__buf_2
XANTENNA__10912__B1 _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1345 net1348 vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__buf_2
XANTENNA__16643__A2 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16811_ _02501_ net104 _02603_ net1712 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[218\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_148_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1356 net1357 vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__clkbuf_2
X_17791_ _08406_ _08407_ _08408_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__and3_2
Xfanout380 _06209_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_2
XANTENNA__13094__S net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_2
X_19530_ clknet_leaf_23_clk game.writer.tracker.next_frame\[125\] net1347 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[125\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11468__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16742_ _02382_ net61 _02582_ net1562 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[170\]
+ sky130_fd_sc_hd__a22o_1
X_13954_ net1052 game.CPU.applesa.ab.check_walls.above.walls\[130\] vssd1 vssd1 vccd1
+ vccd1 _07828_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13862__C1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12905_ game.writer.tracker.frame\[56\] game.writer.tracker.frame\[57\] net1037 vssd1
+ vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__mux2_1
X_19461_ clknet_leaf_39_clk game.writer.tracker.next_frame\[56\] net1352 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[56\] sky130_fd_sc_hd__dfrtp_1
X_16673_ net173 net148 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__nor2_2
X_13885_ net1061 game.CPU.applesa.ab.check_walls.above.walls\[97\] vssd1 vssd1 vccd1
+ vccd1 _07759_ sky130_fd_sc_hd__xor2_1
XANTENNA__12011__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_319_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15603__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18412_ net610 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
X_12836_ game.writer.tracker.frame\[320\] game.writer.tracker.frame\[321\] net1031
+ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__mux2_1
X_15624_ _03483_ net332 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_271_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13614__C1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19392_ clknet_leaf_58_clk _01398_ _00972_ vssd1 vssd1 vccd1 vccd1 game.CPU.bad_collision
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_295_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_335_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09601__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_237_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _01507_ _01542_ _01549_ _01505_ _01574_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__o221a_1
X_18343_ net593 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__inv_2
X_12767_ game.writer.tracker.frame\[116\] game.writer.tracker.frame\[117\] net1026
+ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09833__A1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09833__B2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14506_ _03209_ net1044 net868 game.CPU.apple_location\[4\] _08379_ vssd1 vssd1 vccd1
+ vccd1 _08380_ sky130_fd_sc_hd__o221a_1
XANTENNA__11640__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11718_ net571 _04779_ _05605_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_56_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18274_ net664 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
X_15486_ _08917_ _08931_ _01472_ _01510_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__o211a_1
XANTENNA__11640__B2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15041__C net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12698_ _06560_ _06570_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__nand2_8
XFILLER_0_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13068__S1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17225_ _02541_ net77 _02737_ net1718 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[498\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_13_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14437_ _08307_ _08308_ _08310_ vssd1 vssd1 vccd1 vccd1 _08311_ sky130_fd_sc_hd__or3_1
XANTENNA__17108__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11649_ game.CPU.applesa.ab.check_walls.above.walls\[10\] game.CPU.applesa.ab.apple_possible\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_7_Left_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13393__A1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17156_ _02436_ net59 _02718_ net2034 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[448\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14368_ game.CPU.applesa.ab.absxs.body_x\[117\] net1067 vssd1 vssd1 vccd1 vccd1 _08242_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_268_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19518__Q game.writer.tracker.frame\[113\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12681__B net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16107_ game.CPU.applesa.ab.absxs.body_x\[39\] net461 net443 game.CPU.applesa.ab.absxs.body_y\[38\]
+ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__a22o_1
X_13319_ _06715_ _06717_ _06724_ _06716_ net701 net490 vssd1 vssd1 vccd1 vccd1 _07193_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_326_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17087_ net214 _02393_ net57 _02698_ net1586 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[399\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__10482__A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14299_ _03241_ net1074 _08168_ _08169_ _08172_ vssd1 vssd1 vccd1 vccd1 _08173_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_58_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16038_ game.CPU.applesa.ab.absxs.body_x\[44\] net271 vssd1 vssd1 vccd1 vccd1 _02050_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__14342__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15992__B game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_248_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14889__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13793__A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_271_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18824__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16634__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17989_ net636 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19728_ clknet_leaf_19_clk game.writer.tracker.next_frame\[323\] net1348 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[323\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11459__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12656__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19659_ clknet_leaf_23_clk game.writer.tracker.next_frame\[254\] net1347 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[254\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18974__CLK net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_337_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09412_ net1154 _03449_ _03451_ net1127 _03654_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__a221o_1
XANTENNA__12408__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_259_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13081__A0 _06947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09511__A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ net924 net1268 game.CPU.applesa.ab.absxs.body_y\[90\] net902 vssd1 vssd1
+ vccd1 vccd1 _03586_ sky130_fd_sc_hd__a22o_1
XANTENNA__11760__B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout241_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout339_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09274_ game.CPU.walls.abc.counter vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__inv_2
XFILLER_0_346_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11165__A1_N game.CPU.applesa.ab.absxs.body_y\[50\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1150_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout127_X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16344__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1248_A net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09588__B1 game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17159__B net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_348_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_299_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16063__B net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13179__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_210_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16873__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_A net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11775__X _05663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12811__S net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14151__X _08025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16086__B1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20008__1377 vssd1 vssd1 vccd1 vccd1 net1377 _20008__1377/LO sky130_fd_sc_hd__conb_1
XFILLER_0_356_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__B1 game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ game.CPU.applesa.ab.absxs.body_x\[63\] vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__inv_2
XANTENNA__14311__B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12647__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12112__A game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16389__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_221_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout830_X net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ game.CPU.applesa.ab.absxs.body_x\[29\] net414 net396 game.CPU.applesa.ab.absxs.body_y\[31\]
+ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o221a_1
XANTENNA__16519__A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13642__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09482__A2_N game.CPU.applesa.ab.check_walls.above.walls\[177\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13670_ _07453_ _07454_ _07463_ _07471_ net188 vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__o221a_1
XANTENNA__10673__A2 game.CPU.applesa.ab.absxs.body_x\[115\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11870__A1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10882_ _04780_ _04783_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__or2_1
XFILLER_0_195_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11870__B2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_317_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12621_ _06232_ _06497_ _06233_ _06494_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__or4b_1
XANTENNA__15142__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09815__A1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09815__B2 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ game.writer.updater.commands.cmd_num\[4\] game.writer.updater.commands.cmd_num\[3\]
+ vssd1 vssd1 vccd1 vccd1 _08882_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_182_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12552_ game.CPU.applesa.ab.absxs.body_y\[87\] net364 vssd1 vssd1 vccd1 vccd1 _06429_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16525__Y _02464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ game.CPU.applesa.ab.check_walls.above.walls\[175\] net258 vssd1 vssd1 vccd1
+ vccd1 _05392_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_324_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_310_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15271_ _08812_ _08825_ _08826_ _08815_ _08821_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a32o_1
XFILLER_0_340_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16561__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12483_ game.CPU.applesa.ab.absxs.body_y\[28\] net359 net517 game.CPU.applesa.ab.absxs.body_y\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_163_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17010_ _02501_ net89 _02674_ net1527 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[346\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_297_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13230__X _07104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14222_ game.CPU.applesa.ab.absxs.body_y\[43\] net860 net854 game.CPU.applesa.ab.absxs.body_y\[42\]
+ vssd1 vssd1 vccd1 vccd1 _08096_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_10_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11434_ game.CPU.applesa.ab.check_walls.above.walls\[25\] net771 vssd1 vssd1 vccd1
+ vccd1 _05323_ sky130_fd_sc_hd__xor2_1
XANTENNA__17069__B net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_232_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10389__A1_N net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11398__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14153_ _08015_ _08020_ _08022_ _08026_ vssd1 vssd1 vccd1 vccd1 _08027_ sky130_fd_sc_hd__or4b_4
X_11365_ game.CPU.applesa.ab.check_walls.above.walls\[35\] net763 vssd1 vssd1 vccd1
+ vccd1 _05254_ sky130_fd_sc_hd__xnor2_1
X_13104_ net488 _06977_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__or2_1
X_10316_ _04498_ _04497_ net1843 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__mux2_1
XANTENNA__16864__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18961_ net1201 _00254_ _00632_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_14084_ net942 game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1 vccd1
+ vccd1 _07958_ sky130_fd_sc_hd__xor2_1
X_11296_ _05088_ _05089_ _05092_ _05090_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__or4b_1
XANTENNA__13678__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13817__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13035_ net698 _06876_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__or2_1
X_17912_ net647 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__inv_2
X_10247_ net1166 _04439_ _03362_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__a21oi_1
X_18892_ clknet_leaf_1_clk _01264_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_265_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1120 game.CPU.bodymain1.main.score\[2\] vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_266_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1131 net1132 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__buf_4
X_17843_ game.writer.updater.commands.count\[7\] _08889_ _03165_ vssd1 vssd1 vccd1
+ vccd1 _03169_ sky130_fd_sc_hd__and3_1
Xfanout1142 net1143 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_8_clk_X clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10178_ net1144 _04367_ _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__o21ai_1
Xfanout1153 net1154 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_321_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18997__CLK net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14221__B net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1164 net1165 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_1
XANTENNA__15824__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1175 game.CPU.walls.abc.enable vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__buf_2
Xfanout1186 net1190 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__buf_2
XFILLER_0_206_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17774_ game.CPU.applesa.twoapples.count\[0\] net1163 vssd1 vssd1 vccd1 vccd1 _03125_
+ sky130_fd_sc_hd__and2_1
XANTENNA__15036__C game.CPU.applesa.ab.check_walls.above.walls\[64\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout1197 net1198 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_2
XANTENNA__13835__C1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14986_ net1222 net1250 game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1
+ vccd1 vccd1 _00202_ sky130_fd_sc_hd__and3_1
X_19513_ clknet_leaf_14_clk game.writer.tracker.next_frame\[108\] net1283 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[108\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_178_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09503__B1 game.CPU.applesa.ab.check_walls.above.walls\[50\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16725_ net1953 _02575_ _02577_ net106 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[158\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_282_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13937_ _07800_ _07801_ _07806_ _07810_ vssd1 vssd1 vccd1 vccd1 _07811_ sky130_fd_sc_hd__or4_1
XANTENNA__16429__A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13552__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17041__A2 _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19444_ clknet_leaf_47_clk game.writer.tracker.next_frame\[39\] net1299 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[39\] sky130_fd_sc_hd__dfrtp_1
X_16656_ game.writer.tracker.frame\[120\] _02546_ vssd1 vssd1 vccd1 vccd1 _02547_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_282_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13868_ _06703_ _07545_ _07700_ _07741_ vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_85_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12819_ game.writer.tracker.frame\[326\] game.writer.tracker.frame\[327\] net1026
+ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15607_ game.CPU.applesa.ab.absxs.body_y\[34\] net332 vssd1 vssd1 vccd1 vccd1 _01619_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_186_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19375_ clknet_leaf_9_clk _01381_ _00956_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.snake_head_y\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13799_ net498 _07671_ _07672_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__and3_1
X_16587_ net113 _02387_ _02493_ net728 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__o31a_1
XANTENNA__09806__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09806__B2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12810__A0 game.writer.tracker.frame\[368\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18326_ net599 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
XANTENNA__11613__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15538_ _01540_ _01559_ _01470_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15987__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_332_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19622__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_301_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15469_ game.writer.updater.commands.count\[16\] game.writer.updater.commands.count\[12\]
+ _08892_ _08934_ _01495_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__o311a_1
X_18257_ net644 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_170_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_343_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_343_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17208_ _02525_ net71 net715 vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__o21a_1
XFILLER_0_181_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18188_ net608 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold603 game.CPU.randy.f1.a1.count\[12\] vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11916__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17139_ net158 _02408_ net80 _02714_ net1522 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[435\]
+ sky130_fd_sc_hd__a32o_1
Xhold614 game.writer.tracker.frame\[421\] vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold625 game.CPU.kyle.L1.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 game.writer.tracker.frame\[569\] vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_268_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13118__A1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold647 game.CPU.walls.rand_wall.counter2\[4\] vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 game.writer.tracker.frame\[25\] vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16855__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19772__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09961_ net903 _04186_ _04190_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__nor3_1
Xhold669 game.writer.tracker.frame\[28\] vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16611__B _02480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload26_A clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15508__A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09892_ _03645_ _03647_ _03737_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_168_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17804__A1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09506__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19002__CLK net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout289_A net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17280__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_227_Right_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16134__A1_N game.CPU.applesa.ab.absxs.body_y\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_224_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10104__B2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16339__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13841__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12644__A3 _06515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13315__X _07189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17032__A2 _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1198_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10655__A2 _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12586__B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16058__B _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13054__A0 _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16791__A1 _02470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10387__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout623_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_X net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_270_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09326_ net1096 game.CPU.applesa.ab.absxs.body_x\[81\] vssd1 vssd1 vccd1 vccd1 _03569_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12801__A0 game.writer.tracker.frame\[376\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15897__B net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11080__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ game.CPU.randy.counter1.count1\[8\] vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__inv_2
XFILLER_0_322_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16543__B2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_X net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13357__A1 _06675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13050__X _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09188_ game.CPU.applesa.ab.check_walls.above.walls\[107\] vssd1 vssd1 vccd1 vccd1
+ _03437_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout992_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14306__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14412__A2_N net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17099__A2 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12107__A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13109__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_302_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_268_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16846__A2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11150_ _05034_ _05035_ _05038_ _05039_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__a22o_1
XANTENNA__12317__C1 _06202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_281_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10101_ net1162 _04308_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_73_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11946__A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_79_Left_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11081_ _04963_ _04964_ _04967_ _04968_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__or4_1
X_10032_ _04238_ _04239_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__nor2_1
XANTENNA__09416__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11665__B net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19252__1361 vssd1 vssd1 vccd1 vccd1 _19252__1361/HI net1361 sky130_fd_sc_hd__conb_1
XANTENNA__17271__A2 _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14840_ _08638_ vssd1 vssd1 vccd1 vccd1 _08639_ sky130_fd_sc_hd__inv_2
XFILLER_0_215_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14085__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14771_ net265 _08591_ _08590_ vssd1 vssd1 vccd1 vccd1 _08592_ sky130_fd_sc_hd__o21a_1
XFILLER_0_242_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11983_ game.CPU.applesa.ab.check_walls.above.walls\[180\] net554 vssd1 vssd1 vccd1
+ vccd1 _05870_ sky130_fd_sc_hd__nand2_1
XANTENNA__16249__A net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13832__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13372__S net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_230_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13722_ game.writer.tracker.frame\[195\] net710 net673 game.writer.tracker.frame\[196\]
+ vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__o22a_1
X_16510_ net246 net237 _02325_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_205_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15153__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10934_ game.CPU.applesa.ab.absxs.body_x\[9\] net321 vssd1 vssd1 vccd1 vccd1 _04824_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17490_ net1264 game.CPU.clock1.game_state\[0\] _02782_ _02833_ vssd1 vssd1 vccd1
+ vccd1 _02919_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12496__B net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_88_Left_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09151__A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_292_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16441_ _02283_ net199 _02401_ net239 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__o22a_1
X_13653_ _07525_ _07526_ net483 vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__mux2_1
X_10865_ _03512_ game.CPU.randy.counter1.count1\[3\] _03514_ game.CPU.randy.counter1.count1\[2\]
+ _04743_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__a221o_1
XANTENNA__16782__A1 _02458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19645__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14992__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13596__A1 _07469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_234_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12604_ net1270 net365 net362 game.CPU.applesa.ab.absxs.body_y\[60\] vssd1 vssd1
+ vccd1 vccd1 _06481_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_183_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16372_ net1963 net735 _02352_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[30\]
+ sky130_fd_sc_hd__and3_1
X_19160_ clknet_leaf_3_clk _01281_ _00831_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.counter2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13584_ game.writer.tracker.frame\[339\] net712 net837 game.writer.tracker.frame\[337\]
+ vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10796_ game.CPU.applesa.ab.absxs.body_y\[41\] _04690_ _04728_ game.CPU.applesa.ab.absxs.body_y\[37\]
+ vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__a22o_1
X_15323_ game.CPU.applesa.twomode.counter _08864_ _08865_ _08866_ _08867_ vssd1 vssd1
+ vccd1 vccd1 _08868_ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18111_ net612 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12535_ _06402_ _06403_ _06404_ _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__and4_1
X_19091_ net1178 _00128_ _00762_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[136\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18042_ net659 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__inv_2
X_15254_ _01265_ vssd1 vssd1 vccd1 vccd1 _08813_ sky130_fd_sc_hd__inv_2
XFILLER_0_340_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19795__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12466_ game.CPU.applesa.ab.absxs.body_y\[14\] net520 vssd1 vssd1 vccd1 vccd1 _06343_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_312_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10744__B _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19068__Q game.CPU.applesa.ab.check_walls.above.walls\[113\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14205_ _03268_ net1049 net962 _03335_ _08076_ vssd1 vssd1 vccd1 vccd1 _08079_ sky130_fd_sc_hd__a221o_1
XFILLER_0_340_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11417_ game.CPU.applesa.ab.check_walls.above.walls\[112\] net775 vssd1 vssd1 vccd1
+ vccd1 _05306_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_329_Right_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15185_ _08758_ _08760_ game.CPU.walls.enable_in2 _08754_ vssd1 vssd1 vccd1 vccd1
+ _00085_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_201_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12397_ game.CPU.applesa.ab.absxs.body_y\[93\] net523 vssd1 vssd1 vccd1 vccd1 _06274_
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_97_Left_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14136_ net863 game.CPU.applesa.ab.check_walls.above.walls\[45\] _03405_ net940 vssd1
+ vssd1 vccd1 vccd1 _08010_ sky130_fd_sc_hd__a22o_1
XANTENNA__12571__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11348_ _05236_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19993_ clknet_leaf_45_clk _01417_ net1299 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10582__A1 game.CPU.applesa.ab.absxs.body_x\[115\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12859__A0 _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ net1049 game.CPU.applesa.ab.check_walls.above.walls\[3\] vssd1 vssd1 vccd1
+ vccd1 _07941_ sky130_fd_sc_hd__xor2_1
X_18944_ net1175 _00083_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number_out\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_245_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11279_ _04976_ _04977_ _04978_ _04979_ _05168_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__a221o_2
X_13018_ net506 _06867_ _06868_ _06572_ net680 vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__o221a_1
XANTENNA__09326__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_265_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11575__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20002__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18875_ clknet_leaf_5_clk game.CPU.randy.f1.c1.innerCount\[5\] _00570_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_234_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17262__A2 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17826_ _03150_ _03156_ _03157_ _03146_ game.writer.updater.commands.count\[3\] vssd1
+ vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__a32o_1
XFILLER_0_206_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10885__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19175__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14076__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17757_ game.CPU.applesa.twoapples.count_luck\[2\] _03113_ _03109_ vssd1 vssd1 vccd1
+ vccd1 _03114_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_221_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14969_ game.CPU.walls.rand_wall.logic_enable _08695_ _08742_ _08745_ vssd1 vssd1
+ vccd1 vccd1 _08746_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13282__S net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15063__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17014__A2 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16708_ net174 _02257_ _02328_ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__nor3_1
XFILLER_0_348_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_334_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10637__A2 game.CPU.applesa.ab.absxs.body_x\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17688_ game.CPU.walls.rand_wall.count_luck\[5\] game.CPU.walls.rand_wall.count_luck\[4\]
+ _03068_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__and3_1
XANTENNA__09061__A game.CPU.applesa.ab.absxs.body_y\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19427_ clknet_leaf_41_clk game.writer.tracker.next_frame\[22\] net1330 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_308_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16639_ net131 _02396_ _02516_ _02537_ net1719 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[112\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_202_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16773__A1 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_256_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18374__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_312_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19358_ clknet_leaf_70_clk game.CPU.applesa.twoapples.absxs.next_head\[3\] vssd1
+ vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.x_final\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09111_ net1455 vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20007__1376 vssd1 vssd1 vccd1 vccd1 net1376 _20007__1376/LO sky130_fd_sc_hd__conb_1
XFILLER_0_84_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18309_ net621 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
XFILLER_0_304_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19289_ clknet_leaf_66_clk game.CPU.applesa.ab.absxs.next_head\[7\] vssd1 vssd1 vccd1
+ vccd1 game.CPU.applesa.ab.y_final\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__14407__A game.CPU.applesa.ab.absxs.body_y\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_303_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09042_ game.CPU.applesa.ab.absxs.body_x\[9\] vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__inv_2
XFILLER_0_331_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10654__B _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14000__A2 game.CPU.applesa.ab.check_walls.above.walls\[74\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold400 game.writer.tracker.frame\[114\] vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 game.CPU.randy.f1.a1.count\[7\] vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 game.writer.tracker.frame\[160\] vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_345_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold433 game.writer.tracker.frame\[280\] vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 game.writer.tracker.frame\[501\] vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 game.writer.tracker.frame\[153\] vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 game.writer.tracker.frame\[133\] vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 game.writer.tracker.frame\[490\] vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19355__D game.CPU.applesa.twoapples.absxs.next_head\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18610__Q game.CPU.applesa.ab.absxs.body_y\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold488 game.writer.tracker.frame\[56\] vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout902 net903 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__buf_4
X_09944_ net1114 _04179_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__or2_1
Xhold499 game.writer.tracker.frame\[279\] vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 _03195_ vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__buf_4
XANTENNA__19518__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout924 net925 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__buf_4
XANTENNA__13511__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout935 net937 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_2
Xfanout946 game.CPU.applesa.y\[3\] vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__buf_4
XANTENNA__11485__B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout957 game.CPU.applesa.y\[2\] vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_4
X_09875_ _03552_ _03553_ _03554_ _04019_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__o31a_2
Xfanout968 net972 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10325__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout573_A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 net981 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__buf_4
XANTENNA__13981__A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17253__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_240_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout740_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19668__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout838_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_356_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17005__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16764__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_339_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15701__A game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_354_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18692__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ net1079 _03246_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__nor2_1
XFILLER_0_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16516__B net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13673__S1 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ net1142 _03306_ _03307_ net1149 _03550_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_354_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10581_ net1080 _04663_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__nor2_2
XFILLER_0_180_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12320_ _06142_ _06143_ _06144_ _06136_ _06135_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__o32a_1
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10800__A2 _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19048__CLK net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ net804 net549 vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16532__A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_309_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11202_ _03249_ net320 vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__xnor2_1
X_12182_ game.CPU.applesa.ab.check_walls.above.walls\[61\] net550 vssd1 vssd1 vccd1
+ vccd1 _06068_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_151_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10564__A1 game.CPU.applesa.ab.absxs.body_x\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16251__B net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11133_ game.CPU.applesa.ab.absxs.body_x\[69\] net322 vssd1 vssd1 vccd1 vccd1 _05023_
+ sky130_fd_sc_hd__or2_1
XANTENNA__15148__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16295__A3 _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16990_ _02473_ net86 net715 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__o21a_1
XFILLER_0_275_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13502__A1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09146__A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ _03281_ net326 vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__xnor2_1
X_15941_ net821 net439 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__nor2_1
XANTENNA__11395__B net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _04219_ _04222_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_262_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17244__A2 _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18660_ clknet_leaf_60_clk _01077_ _00397_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[78\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_250_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15872_ _03349_ net333 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__xnor2_1
X_17611_ game.CPU.kyle.L1.cnt_20ms\[9\] game.CPU.kyle.L1.cnt_20ms\[8\] _03020_ vssd1
+ vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__and3_1
X_14823_ game.CPU.randy.counter1.count\[16\] _08626_ vssd1 vssd1 vccd1 vccd1 _08629_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_263_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18591_ clknet_leaf_50_clk _01011_ _00328_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[64\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_240_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13361__S0 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17542_ game.CPU.modea.Qa\[0\] _02845_ _02856_ game.CPU.kyle.L1.row_2\[72\] _02968_
+ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11816__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11966_ _05731_ _05752_ _05770_ _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__or4_1
X_14754_ game.CPU.randy.counter1.count1\[17\] _08575_ vssd1 vssd1 vccd1 vccd1 _08577_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_230_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14304__A2_N net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13705_ _07577_ _07578_ net487 vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__mux2_1
X_10917_ net411 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.next_head\[2\] sky130_fd_sc_hd__inv_2
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17473_ _03198_ _02786_ _02787_ _02802_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__o22a_1
X_14685_ game.CPU.randy.counter1.count1\[11\] _08491_ _08502_ game.CPU.randy.counter1.count1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _08524_ sky130_fd_sc_hd__o22ai_1
XANTENNA__16755__A1 _02404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11897_ net573 _05409_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__nor2_1
XFILLER_0_357_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19212_ net1167 _00024_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_possible\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13636_ game.writer.tracker.frame\[23\] net711 net674 game.writer.tracker.frame\[24\]
+ _07509_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__o221a_1
X_16424_ net163 _02389_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__and2_2
XFILLER_0_345_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10848_ _03503_ game.CPU.randy.counter1.count1\[10\] _03504_ game.CPU.randy.counter1.count1\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16426__B _02310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19143_ net1184 _00185_ _00814_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[188\]
+ sky130_fd_sc_hd__dfrtp_1
X_16355_ _02247_ net235 _02283_ _02339_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__o31a_4
X_13567_ _07439_ _07440_ net500 vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__mux2_1
XANTENNA__16507__B2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10779_ _03306_ net327 vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__nor2_1
X_12518_ game.CPU.applesa.ab.absxs.body_x\[69\] net379 vssd1 vssd1 vccd1 vccd1 _06395_
+ sky130_fd_sc_hd__and2_1
X_15306_ _08853_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_325_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_298_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16286_ net239 _02227_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19074_ net1186 _00109_ _00745_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[119\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13498_ _07370_ _07371_ net514 vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__mux2_1
XANTENNA__17180__A1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_251_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_288_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18025_ net662 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__inv_2
XFILLER_0_301_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15237_ net1415 _03490_ net1282 vssd1 vssd1 vccd1 vccd1 _08799_ sky130_fd_sc_hd__o21ai_4
X_12449_ _03273_ game.CPU.applesa.twoapples.absxs.next_head\[0\] vssd1 vssd1 vccd1
+ vccd1 _06326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_313_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_288_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15168_ net1227 net1254 game.CPU.walls.rand_wall.y_final\[0\] vssd1 vssd1 vccd1 vccd1
+ _00232_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14119_ _07984_ _07985_ _07989_ _07990_ vssd1 vssd1 vccd1 vccd1 _07993_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_35_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15058__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19976_ clknet_leaf_41_clk game.writer.tracker.next_frame\[571\] net1330 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[571\] sky130_fd_sc_hd__dfrtp_1
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_2
X_15099_ net1203 net1229 game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1
+ vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14297__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18927_ clknet_leaf_4_clk net1408 _00611_ vssd1 vssd1 vccd1 vccd1 game.CPU.right_button.eD1.Q2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_293_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18565__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14897__A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_340_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_307_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17235__A2 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19810__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09660_ _03898_ _03899_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__or3_4
X_18858_ clknet_leaf_1_clk _01249_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_253_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17809_ _08883_ _08934_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09591_ net923 game.CPU.applesa.ab.check_walls.above.walls\[18\] game.CPU.applesa.ab.check_walls.above.walls\[20\]
+ net894 _03833_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__o221a_1
XANTENNA__10489__X _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18789_ clknet_leaf_4_clk _01204_ _00526_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13306__A net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11807__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12210__A game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19960__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout154_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15521__A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_176_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_336_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_351_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_336_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11035__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout321_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10665__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1063_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout419_A net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10243__B1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17171__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09025_ game.CPU.applesa.ab.absxs.body_x\[43\] vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout207_X net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_304_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1328_A net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19340__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold230 game.writer.tracker.frame\[478\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 game.CPU.randy.f1.c1.count\[10\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 game.writer.tracker.frame\[507\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout690_A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10671__Y _04702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16071__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 game.writer.tracker.frame\[222\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_265_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout788_A game.CPU.applesa.ab.check_walls.above.walls\[159\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18908__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 game.writer.tracker.frame\[124\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 game.writer.tracker.frame\[141\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_348_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold296 game.writer.tracker.frame\[46\] vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_217_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout710 net712 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__buf_4
XANTENNA__15485__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14288__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_X clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout721 net726 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout732 net733 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_187_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09927_ _04150_ _04166_ net1261 vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__a21bo_1
Xfanout743 _04451_ vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout955_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout754 _04159_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__buf_6
XANTENNA__18279__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19490__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout765 net767 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_129_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17226__A2 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout776 game.CPU.applesa.ab.apple_possible\[0\] vssd1 vssd1 vccd1 vccd1 net776
+ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_304_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13591__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09858_ net1112 game.CPU.applesa.ab.absxs.body_x\[44\] vssd1 vssd1 vccd1 vccd1 _04101_
+ sky130_fd_sc_hd__xor2_1
Xfanout787 game.CPU.applesa.ab.check_walls.above.walls\[166\] vssd1 vssd1 vccd1 vccd1
+ net787 sky130_fd_sc_hd__clkbuf_4
X_20047_ game.CPU.applesa.ab.good_collision vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
Xfanout798 game.CPU.applesa.ab.check_walls.above.walls\[117\] vssd1 vssd1 vccd1 vccd1
+ net798 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout67_A _02393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11943__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09789_ _04026_ _04027_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16985__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_clk_X clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16985__B2 game.writer.tracker.frame\[329\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11820_ net826 net393 net308 game.CPU.applesa.ab.check_walls.above.walls\[29\] _05707_
+ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__a221o_1
XFILLER_0_197_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12120__A game.CPU.applesa.ab.check_walls.above.walls\[172\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_202_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_276_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ net748 _05385_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16737__A1 _02369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_233_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13503__X _07377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_218_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14973__C game.CPU.applesa.ab.check_walls.above.walls\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10702_ game.CPU.applesa.ab.absxs.body_y\[76\] _04623_ _04624_ game.CPU.applesa.ab.absxs.body_y\[72\]
+ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__a22o_1
X_14470_ _08336_ _08343_ _08342_ _08341_ vssd1 vssd1 vccd1 vccd1 _08344_ sky130_fd_sc_hd__or4b_1
XFILLER_0_138_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11682_ net778 _05570_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__xor2_1
X_13421_ _06600_ _06994_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__or2_1
X_10633_ game.CPU.applesa.ab.absxs.body_x\[56\] net328 _04684_ net935 vssd1 vssd1
+ vccd1 vccd1 _01119_ sky130_fd_sc_hd__a22o_1
XANTENNA__15150__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14047__A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16140_ net1267 net356 net352 _03236_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__o2bb2a_1
X_13352_ _06644_ _06655_ _06656_ _06657_ net509 net701 vssd1 vssd1 vccd1 vccd1 _07226_
+ sky130_fd_sc_hd__mux4_1
X_10564_ game.CPU.applesa.ab.absxs.body_x\[15\] _04653_ _04654_ game.CPU.applesa.ab.absxs.body_x\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__a22o_1
XANTENNA__17162__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12303_ net821 net419 vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__xnor2_1
X_16071_ _03232_ net465 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__nand2_1
X_13283_ _07152_ _07155_ net683 vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_350_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16262__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10495_ net1120 net1124 net1122 net1118 vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__or4bb_1
X_15022_ net1222 net1256 game.CPU.applesa.ab.check_walls.above.walls\[50\] vssd1 vssd1
+ vccd1 vccd1 _00241_ sky130_fd_sc_hd__and3_1
X_12234_ game.CPU.applesa.ab.check_walls.above.walls\[71\] net423 vssd1 vssd1 vccd1
+ vccd1 _06120_ sky130_fd_sc_hd__nand2_1
XANTENNA__11677__Y _05566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10537__A1 game.CPU.applesa.ab.absxs.body_x\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_287_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18588__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11734__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19830_ clknet_leaf_38_clk game.writer.tracker.next_frame\[425\] net1325 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[425\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19833__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ game.CPU.applesa.ab.check_walls.above.walls\[156\] net552 vssd1 vssd1 vccd1
+ vccd1 _06052_ sky130_fd_sc_hd__nand2_1
XFILLER_0_258_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_229_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14279__A2 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11116_ _04996_ _05000_ _05004_ _05005_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__or4_1
X_19761_ clknet_leaf_30_clk game.writer.tracker.next_frame\[356\] net1313 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[356\] sky130_fd_sc_hd__dfrtp_1
X_16973_ net1515 _02662_ _02442_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[321\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_275_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17805__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12096_ net802 net296 net290 net803 vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_263_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11693__X _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18712_ clknet_leaf_60_clk _01129_ _00449_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[74\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13582__S0 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17217__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ _03329_ net403 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__xnor2_1
X_15924_ game.CPU.applesa.ab.check_walls.above.walls\[130\] net346 vssd1 vssd1 vccd1
+ vccd1 _01936_ sky130_fd_sc_hd__or2_1
X_19692_ clknet_leaf_26_clk game.writer.tracker.next_frame\[287\] net1313 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[287\] sky130_fd_sc_hd__dfrtp_1
X_20006__1375 vssd1 vssd1 vccd1 vccd1 net1375 _20006__1375/LO sky130_fd_sc_hd__conb_1
XFILLER_0_204_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16425__B1 _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19983__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18643_ clknet_leaf_53_clk _01060_ _00380_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[45\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_30_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _03260_ game.CPU.walls.rand_wall.abduyd.next_wall\[3\] net340 _03325_ vssd1
+ vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a22o_1
XANTENNA__15779__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14806_ game.CPU.randy.counter1.count\[10\] _08616_ net138 vssd1 vssd1 vccd1 vccd1
+ _08618_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_318_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18574_ clknet_leaf_62_clk _00994_ _00311_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_15786_ _03331_ net440 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__nand2_1
X_12998_ game.writer.tracker.frame\[526\] game.writer.tracker.frame\[527\] net1006
+ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10469__B net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17525_ _02845_ _02950_ _02949_ _02855_ _02850_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_129_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16728__A1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19213__CLK net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14737_ _03502_ _08563_ vssd1 vssd1 vccd1 vccd1 _08566_ sky130_fd_sc_hd__nand2_1
X_11949_ net749 _05302_ _05306_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_71_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_290_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17456_ _02787_ _02792_ net1117 _02785_ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_253_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14668_ _04348_ net266 game.CPU.randy.counter1.count1\[6\] vssd1 vssd1 vccd1 vccd1
+ _08507_ sky130_fd_sc_hd__o21a_1
XANTENNA__14203__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16407_ net196 _02376_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__nor2_2
X_13619_ game.writer.tracker.frame\[285\] game.writer.tracker.frame\[287\] game.writer.tracker.frame\[288\]
+ game.writer.tracker.frame\[286\] net976 net1012 vssd1 vssd1 vccd1 vccd1 _07493_
+ sky130_fd_sc_hd__mux4_1
X_17387_ _03217_ game.CPU.kyle.L1.nextState\[2\] vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__and2_1
XFILLER_0_333_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14599_ game.CPU.clock1.counter\[3\] _08455_ game.CPU.clock1.counter\[4\] vssd1 vssd1
+ vccd1 vccd1 _08457_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_306_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19363__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19126_ net1183 _00167_ _00797_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[171\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13962__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16338_ net238 _02244_ net236 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__or3_4
XFILLER_0_109_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17153__A1 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13962__B2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16443__Y _02404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19057_ net1191 _00091_ _00728_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[102\]
+ sky130_fd_sc_hd__dfrtp_2
X_16269_ net162 _02271_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__nor2_4
XANTENNA__16900__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_329_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_313_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_285_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18008_ net616 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__inv_2
XANTENNA__09918__B1 _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10528__A1 game.CPU.applesa.ab.absxs.body_x\[54\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10932__B net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_239_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_273_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19959_ clknet_leaf_44_clk game.writer.tracker.next_frame\[554\] net1303 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[554\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18099__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09712_ net916 game.CPU.applesa.ab.absxs.body_x\[21\] _03317_ net1158 vssd1 vssd1
+ vccd1 vccd1 _03955_ sky130_fd_sc_hd__a22o_1
XANTENNA__17208__A2 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13573__S0 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_241_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09643_ _03883_ _03884_ _03885_ _03882_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__a211o_1
XFILLER_0_207_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16967__A1 _02429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout271_A net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10700__A1 game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_A game.CPU.applesa.twoapples.absxs.next_head\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10700__B2 game.CPU.applesa.ab.absxs.body_y\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_96_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09574_ net1110 game.CPU.applesa.ab.check_walls.above.walls\[40\] vssd1 vssd1 vccd1
+ vccd1 _03817_ sky130_fd_sc_hd__xor2_1
XFILLER_0_210_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_353_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_328_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_309_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16719__B2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout157_X net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_60_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19706__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16066__B _08429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout703_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_X net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13953__A1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17144__A1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13953__B2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10767__B2 game.CPU.applesa.ab.absxs.body_y\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11964__B1 _05819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18730__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19856__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12814__S net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14154__X _08028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16082__A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09008_ game.CPU.applesa.ab.absxs.body_x\[111\] vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__inv_2
X_10280_ _04256_ _04436_ _04440_ _04471_ _04472_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.good_spot_next
+ sky130_fd_sc_hd__o32a_4
XTAP_TAPCELL_ROW_306_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14314__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17906__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15129__C game.CPU.applesa.ab.check_walls.above.walls\[157\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16655__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18880__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_X net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_4
Xfanout551 net555 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_2
XFILLER_0_272_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout562 _04629_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_217_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13970_ net867 net810 _03426_ net939 _07843_ vssd1 vssd1 vccd1 vccd1 _07844_ sky130_fd_sc_hd__o221a_1
Xfanout573 net575 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_13_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout584 net585 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__buf_2
Xfanout595 net598 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_2
X_12921_ net212 _06695_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__and2_2
XFILLER_0_232_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15145__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11673__B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16958__A1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19236__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_224_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15713__X _01725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15640_ _03266_ net269 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__xnor2_1
X_12852_ game.writer.tracker.frame\[266\] game.writer.tracker.frame\[267\] net996
+ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16528__Y _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14984__B net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_240_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11803_ game.CPU.applesa.ab.check_walls.above.walls\[61\] net308 vssd1 vssd1 vccd1
+ vccd1 _05691_ sky130_fd_sc_hd__nand2_1
X_12783_ game.writer.tracker.frame\[94\] game.writer.tracker.frame\[95\] net1017 vssd1
+ vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__mux2_1
XANTENNA__12444__A1 game.CPU.applesa.ab.absxs.body_y\[106\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15571_ net1427 net1420 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_28_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12444__B2 game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_346_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17310_ net130 _02535_ net1948 net724 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[561\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15161__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14522_ _08395_ vssd1 vssd1 vccd1 vccd1 _08396_ sky130_fd_sc_hd__inv_2
X_11734_ net749 _05478_ net392 game.CPU.applesa.ab.check_walls.above.walls\[108\]
+ _05620_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__a221o_1
XANTENNA__19386__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18290_ net618 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16186__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17241_ _02551_ net79 _02741_ net1745 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[510\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_202_Left_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14453_ _03251_ net1067 net858 game.CPU.applesa.ab.absxs.body_y\[15\] vssd1 vssd1
+ vccd1 vccd1 _08327_ sky130_fd_sc_hd__o22a_1
X_11665_ game.CPU.applesa.ab.check_walls.above.walls\[121\] net769 vssd1 vssd1 vccd1
+ vccd1 _05554_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_315_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_289_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13404_ _07274_ _07277_ net225 vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__mux2_1
XANTENNA__13944__A1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10616_ game.CPU.applesa.ab.absxs.body_x\[73\] _04675_ _04676_ game.CPU.applesa.ab.absxs.body_x\[69\]
+ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__a22o_1
X_17172_ _02468_ net71 net715 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__o21a_1
XANTENNA__13944__B2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14384_ _08251_ _08255_ _08256_ _08257_ vssd1 vssd1 vccd1 vccd1 _08258_ sky130_fd_sc_hd__and4_1
XANTENNA__17135__A1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11596_ game.CPU.applesa.ab.check_walls.above.walls\[109\] net315 vssd1 vssd1 vccd1
+ vccd1 _05485_ sky130_fd_sc_hd__or2_1
XANTENNA__17135__B2 game.writer.tracker.frame\[432\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10758__A1 game.CPU.applesa.ab.absxs.body_y\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12009__B net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13335_ net239 _07203_ _07208_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__and3_1
X_16123_ game.CPU.applesa.ab.absxs.body_x\[54\] net467 net334 _03306_ vssd1 vssd1
+ vccd1 vccd1 _02135_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10547_ net1117 _03198_ net1121 _04607_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__or4_1
XFILLER_0_106_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_268_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15697__A1 game.CPU.applesa.ab.absxs.body_x\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_267_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15697__B2 game.CPU.applesa.ab.absxs.body_y\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13266_ game.writer.tracker.frame\[482\] game.writer.tracker.frame\[483\] net1011
+ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__mux2_1
XANTENNA__11848__B net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16054_ game.CPU.applesa.ab.absxs.body_x\[102\] net469 net440 game.CPU.applesa.ab.absxs.body_y\[102\]
+ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__a22o_1
X_10478_ game.CPU.applesa.ab.absxs.body_x\[92\] _04601_ _04605_ net929 vssd1 vssd1
+ vccd1 vccd1 _01195_ sky130_fd_sc_hd__a22o_1
XANTENNA__19076__Q game.CPU.applesa.ab.check_walls.above.walls\[121\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14224__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_295_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15005_ net1221 net1249 game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1 vssd1
+ vccd1 vccd1 _00223_ sky130_fd_sc_hd__and3_1
X_12217_ _06013_ _06102_ _06015_ _06014_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_283_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13197_ net231 _07070_ _07065_ net279 vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_90_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12025__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15039__C game.CPU.applesa.ab.check_walls.above.walls\[67\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19813_ clknet_leaf_37_clk game.writer.tracker.next_frame\[408\] net1349 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[408\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_236_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17094__Y _02700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12148_ _05458_ _05459_ _05460_ _05461_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_211_Left_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16110__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_324_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19744_ clknet_leaf_24_clk game.writer.tracker.next_frame\[339\] net1340 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[339\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14121__B2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16661__A3 _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16956_ net155 _02413_ net86 net729 vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__o31a_1
XFILLER_0_208_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ net809 net289 vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__xor2_1
XANTENNA__12312__X _06198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12132__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15907_ game.CPU.applesa.ab.absxs.body_y\[56\] net452 vssd1 vssd1 vccd1 vccd1 _01919_
+ sky130_fd_sc_hd__xnor2_1
X_19675_ clknet_leaf_32_clk game.writer.tracker.next_frame\[270\] net1285 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[270\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11486__A2 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16887_ _02240_ _02634_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18626_ clknet_leaf_16_clk _01043_ _00363_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_0_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _03388_ net468 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__nand2_1
XANTENNA__18603__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19729__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14424__A2 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_304_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18557_ clknet_leaf_1_clk _00013_ _00294_ vssd1 vssd1 vccd1 vccd1 game.CPU.speed1.Qa\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13632__B1 net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15769_ _01774_ _01776_ _01779_ _01780_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__or4_1
XFILLER_0_63_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09300__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17508_ _02775_ _02842_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__nor2_1
XANTENNA__09300__B2 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09290_ net1156 net810 vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__nand2_1
X_18488_ net583 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16177__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10927__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17439_ _02836_ _02862_ _02864_ _02868_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__or4_1
XANTENNA_14 _02998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18753__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19879__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12982__X _06856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _07032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18382__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_36 _08359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13396__C1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 _08416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11104__A game.CPU.applesa.ab.absxs.body_x\[35\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17126__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload56_A clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19109_ net1181 _00148_ _00780_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[154\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11410__A2 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout117_A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13148__C1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09509__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13699__B1 _07569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14360__A1 net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14360__B2 net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_262_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16637__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13465__S net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_A _06596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14112__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14112__B2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12123__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13320__C1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_301_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17062__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09626_ net1130 game.CPU.applesa.ab.absxs.body_y\[19\] vssd1 vssd1 vccd1 vccd1 _03869_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_179_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_329_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_250_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09531__X _03774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09557_ net913 game.CPU.applesa.ab.absxs.body_x\[60\] net1270 net908 vssd1 vssd1
+ vccd1 vccd1 _03800_ sky130_fd_sc_hd__o22a_1
XFILLER_0_195_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout441_X net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_X net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_328_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10437__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_273_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09488_ net1082 game.CPU.applesa.ab.check_walls.above.walls\[187\] vssd1 vssd1 vccd1
+ vccd1 _03731_ sky130_fd_sc_hd__xor2_1
XANTENNA__16168__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_195_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_230_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11450_ net565 _05338_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_137_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_312_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17117__A1 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20005__1374 vssd1 vssd1 vccd1 vccd1 net1374 _20005__1374/LO sky130_fd_sc_hd__conb_1
X_10401_ net1260 game.CPU.randy.f1.state\[4\] _04360_ _04547_ vssd1 vssd1 vccd1 vccd1
+ _04551_ sky130_fd_sc_hd__or4b_1
XFILLER_0_190_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11381_ game.CPU.applesa.ab.check_walls.above.walls\[176\] net775 vssd1 vssd1 vccd1
+ vccd1 _05270_ sky130_fd_sc_hd__xor2_1
XFILLER_0_104_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14325__A game.CPU.applesa.ab.absxs.body_y\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_277_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ game.writer.tracker.frame\[174\] game.writer.tracker.frame\[175\] net991
+ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_249_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10332_ _04487_ _04492_ _04507_ net739 net1926 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__a32o_1
XANTENNA__09419__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14044__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10572__B net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Left_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13051_ game.writer.tracker.frame\[250\] game.writer.tracker.frame\[251\] net1031
+ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_284_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10263_ net1173 _04394_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16540__A net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ game.CPU.applesa.ab.check_walls.above.walls\[164\] net552 vssd1 vssd1 vccd1
+ vccd1 _05889_ sky130_fd_sc_hd__or2_1
XANTENNA__11165__B2 game.CPU.applesa.ab.absxs.body_x\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_226_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1302 net1307 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13883__B game.CPU.applesa.ab.check_walls.above.walls\[98\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10194_ net1108 _04381_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__nand2_1
Xfanout1313 net1314 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__clkbuf_4
Xfanout1324 net1325 vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__clkbuf_4
Xfanout1335 net1337 vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__clkbuf_4
X_16810_ net150 _02498_ net104 _02603_ net1710 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[217\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__15156__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11684__A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1346 net1347 vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13537__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1357 net1358 vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16643__A3 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_233_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14060__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17790_ _08813_ _08837_ _03133_ _08812_ vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__o211a_1
XFILLER_0_260_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18626__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout370 net374 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_4
XANTENNA__13311__C1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout381 net385 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_260_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16741_ _02378_ net101 _02582_ net1705 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[169\]
+ sky130_fd_sc_hd__a22o_1
Xfanout392 net395 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_4
X_13953_ net1069 _03447_ _03450_ net947 _07822_ vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__a221o_1
XANTENNA__13862__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14995__A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18467__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11971__X _05858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19460_ clknet_leaf_39_clk game.writer.tracker.next_frame\[55\] net1352 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[55\] sky130_fd_sc_hd__dfrtp_1
X_12904_ _06774_ _06775_ _06777_ _06776_ net495 net685 vssd1 vssd1 vccd1 vccd1 _06778_
+ sky130_fd_sc_hd__mux4_1
X_16672_ net134 _02257_ _02357_ net718 vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__o31a_1
XANTENNA__13912__A2_N game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13884_ net1046 game.CPU.applesa.ab.check_walls.above.walls\[99\] vssd1 vssd1 vccd1
+ vccd1 _07758_ sky130_fd_sc_hd__xor2_1
XANTENNA__08993__A game.CPU.applesa.ab.absxs.body_x\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_213_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16800__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09441__X _03684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18411_ net610 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__inv_2
X_15623_ game.CPU.applesa.ab.absxs.body_x\[70\] net467 vssd1 vssd1 vccd1 vccd1 _01635_
+ sky130_fd_sc_hd__xnor2_1
X_12835_ game.writer.tracker.frame\[316\] game.writer.tracker.frame\[317\] net1032
+ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18776__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19391_ clknet_leaf_9_clk _01397_ _00971_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.snake_head_x\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_295_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_271_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10428__B1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18342_ net595 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _06551_ _06585_ _01508_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__or3_1
XANTENNA__09601__B game.CPU.applesa.ab.absxs.body_x\[73\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12766_ game.writer.tracker.frame\[120\] game.writer.tracker.frame\[121\] net1030
+ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_237_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14505_ _03210_ net1060 net856 game.CPU.apple_location\[7\] vssd1 vssd1 vccd1 vccd1
+ _08379_ sky130_fd_sc_hd__o22a_1
XFILLER_0_327_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18273_ net662 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
X_11717_ game.CPU.applesa.ab.apple_possible\[4\] net759 net571 game.CPU.applesa.ab.apple_possible\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__a31o_1
X_12697_ _06560_ _06570_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__and2_4
X_15485_ net993 _01506_ _01508_ net1076 _01509_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__o221a_1
XFILLER_0_126_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16715__A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17224_ _02539_ _02720_ net727 vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__o21a_1
XANTENNA__13917__A1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13917__B2 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14436_ _03279_ net1054 net959 _03350_ _08309_ vssd1 vssd1 vccd1 vccd1 _08310_ sky130_fd_sc_hd__a221o_1
X_11648_ game.CPU.applesa.ab.check_walls.above.walls\[8\] net778 vssd1 vssd1 vccd1
+ vccd1 _05537_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_13_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16434__B net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17155_ _02435_ net58 _02718_ net1602 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[447\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_181_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14367_ game.CPU.applesa.ab.absxs.body_x\[119\] net1050 vssd1 vssd1 vccd1 vccd1 _08241_
+ sky130_fd_sc_hd__xor2_1
X_11579_ net563 _05459_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__or2_1
XANTENNA__14235__A game.CPU.applesa.ab.absxs.body_y\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16106_ _02112_ _02113_ _02116_ _02117_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__or4_2
X_13318_ net686 _06723_ _07191_ net228 vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_326_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17086_ _02257_ _02479_ net71 net735 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__o31a_1
X_14298_ game.CPU.applesa.ab.absxs.body_y\[52\] net871 _08165_ _08166_ _08171_ vssd1
+ vssd1 vccd1 vccd1 _08172_ sky130_fd_sc_hd__a2111o_1
XANTENNA__16721__Y _02576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09349__A1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19401__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_208_Right_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_311_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16037_ _02045_ _02046_ _02047_ _02048_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__or4_1
XANTENNA__09349__B2 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13249_ game.writer.tracker.frame\[468\] game.writer.tracker.frame\[469\] net1014
+ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_255_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_248_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_296_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19534__Q game.writer.tracker.frame\[129\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13528__S0 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16634__A3 _02391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17988_ net634 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12105__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19551__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19727_ clknet_leaf_19_clk game.writer.tracker.next_frame\[322\] net1348 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[322\] sky130_fd_sc_hd__dfrtp_1
X_16939_ net148 _02530_ net86 net713 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__o31a_1
XANTENNA__11459__A2 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12202__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_108_Left_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_315_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11881__X _05769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19658_ clknet_leaf_23_clk game.writer.tracker.next_frame\[253\] net1347 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[253\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10003__A net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_337_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09411_ net1108 game.CPU.applesa.ab.check_walls.above.walls\[128\] vssd1 vssd1 vccd1
+ vccd1 _03654_ sky130_fd_sc_hd__xor2_1
X_18609_ clknet_leaf_70_clk _01026_ _00346_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[91\]
+ sky130_fd_sc_hd__dfrtp_4
X_19589_ clknet_leaf_36_clk game.writer.tracker.next_frame\[184\] net1354 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[184\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13605__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12408__B2 game.CPU.applesa.ab.absxs.body_y\[52\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_17_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_259_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09342_ net924 net1268 _03326_ net1136 vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_121_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13700__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09273_ game.CPU.clock1.counter\[21\] vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__inv_2
XANTENNA__16184__X _02196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16625__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout234_A _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14030__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16344__B _02258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_117_Left_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19358__D game.CPU.applesa.twoapples.absxs.next_head\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09588__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout401_A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_210_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_348_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09239__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19081__CLK net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_302_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_307_Left_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_247_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1310_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16360__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18649__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__B2 game.CPU.applesa.ab.absxs.body_x\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout770_A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13195__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A _03374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16086__B2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__B2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08988_ game.CPU.applesa.ab.absxs.body_x\[71\] vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__inv_2
XANTENNA__10370__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Left_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18287__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12112__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12631__A1_N game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_199_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10950_ _03248_ net323 net411 game.CPU.applesa.ab.absxs.body_x\[30\] vssd1 vssd1
+ vccd1 vccd1 _04840_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_221_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16389__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_316_Left_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09609_ net1149 game.CPU.applesa.ab.absxs.body_y\[117\] vssd1 vssd1 vccd1 vccd1 _03852_
+ sky130_fd_sc_hd__xor2_1
X_10881_ game.CPU.applesa.ab.apple_possible\[6\] _04779_ vssd1 vssd1 vccd1 vccd1 _04783_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11870__A2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12620_ game.CPU.applesa.ab.absxs.body_x\[79\] net531 net526 game.CPU.applesa.ab.absxs.body_y\[77\]
+ _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__a221o_1
XFILLER_0_344_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_316_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12551_ game.CPU.applesa.ab.absxs.body_y\[11\] net366 vssd1 vssd1 vccd1 vccd1 _06428_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_309_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_241_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14981__C game.CPU.applesa.ab.check_walls.above.walls\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11502_ net785 net250 _05380_ _05389_ _05390_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__o2111a_1
XANTENNA__10830__A0 net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_135_Left_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12482_ game.CPU.applesa.ab.absxs.body_x\[29\] net375 net369 _03315_ vssd1 vssd1
+ vccd1 vccd1 _06359_ sky130_fd_sc_hd__o22a_1
X_15270_ _08819_ _08820_ _08824_ vssd1 vssd1 vccd1 vccd1 _08826_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16561__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09579__A1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19424__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11433_ _05321_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__inv_2
X_14221_ game.CPU.applesa.ab.absxs.body_y\[41\] net961 vssd1 vssd1 vccd1 vccd1 _08095_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_10_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09579__B2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_269_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14055__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14572__B2 _00039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_232_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11386__A1 game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_312_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14152_ _07799_ _08023_ _08024_ _08025_ vssd1 vssd1 vccd1 vccd1 _08026_ sky130_fd_sc_hd__and4_1
XANTENNA__09149__A game.CPU.applesa.ab.check_walls.above.walls\[35\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_325_Left_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11364_ game.CPU.applesa.ab.check_walls.above.walls\[35\] net763 vssd1 vssd1 vccd1
+ vccd1 _05253_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15588__A1_N net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13103_ _06930_ _06933_ net682 vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__mux2_1
X_10315_ game.CPU.randy.f1.a1.count\[14\] _04487_ _04495_ vssd1 vssd1 vccd1 vccd1
+ _04498_ sky130_fd_sc_hd__and3_1
XANTENNA__11966__X _05854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18960_ net1201 _00243_ _00631_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_14083_ net1063 game.CPU.applesa.ab.check_walls.above.walls\[89\] vssd1 vssd1 vccd1
+ vccd1 _07957_ sky130_fd_sc_hd__xor2_1
XANTENNA__16270__A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11295_ _04913_ _04914_ _05183_ _05184_ _04844_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__o41a_2
XFILLER_0_265_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13034_ _06874_ _06889_ net698 vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__mux2_1
X_17911_ net647 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__inv_2
X_10246_ _04434_ _04438_ _04428_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_265_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18891_ clknet_leaf_2_clk _01263_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__19840__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1110 net1113 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__buf_4
XANTENNA__09751__A1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1121 net1123 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_2
X_17842_ game.writer.updater.commands.count\[8\] _03166_ _03168_ net182 _03155_ vssd1
+ vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__o221a_1
Xfanout1132 net1133 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_266_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09751__B2 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ net1153 _04369_ _04368_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_206_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1143 game.CPU.applesa.ab.snake_head_y\[2\] vssd1 vssd1 vccd1 vccd1 net1143
+ sky130_fd_sc_hd__buf_4
Xfanout1154 net1157 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_321_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1165 game.CPU.applesa.enablea2 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__buf_2
Xfanout1176 game.CPU.walls.abc.enable vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_4
X_17773_ _03109_ _03123_ _03124_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__and3_1
Xfanout1187 net1188 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__buf_2
X_14985_ net1224 net1251 game.CPU.applesa.ab.check_walls.above.walls\[13\] vssd1 vssd1
+ vccd1 vccd1 _00201_ sky130_fd_sc_hd__and3_1
Xfanout1198 net1202 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17026__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_233_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19512_ clknet_leaf_14_clk game.writer.tracker.next_frame\[107\] net1283 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[107\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09503__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16724_ _02257_ _02430_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__nor2_2
XANTENNA__15614__A game.CPU.applesa.ab.check_walls.above.walls\[83\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09503__B2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_334_Left_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13936_ net1072 _03396_ _03398_ net1046 _07809_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__a221o_1
XFILLER_0_214_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_282_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19443_ clknet_leaf_47_clk game.writer.tracker.next_frame\[38\] net1299 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[38\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11861__B net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16655_ net114 _02545_ net730 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__o21a_1
XFILLER_0_186_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15588__B1 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13867_ net184 net174 _07740_ net162 vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10664__A3 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_347_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15606_ _01609_ _01614_ _01615_ _01617_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__or4_2
X_12818_ game.writer.tracker.frame\[322\] game.writer.tracker.frame\[323\] net1030
+ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_215_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19374_ clknet_leaf_71_clk _01380_ _00955_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17329__A1 _02275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16586_ net197 _02387_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__nor2_1
XANTENNA__15052__C game.CPU.applesa.ab.check_walls.above.walls\[80\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ game.writer.tracker.frame\[386\] net843 net673 game.writer.tracker.frame\[388\]
+ vssd1 vssd1 vccd1 vccd1 _07672_ sky130_fd_sc_hd__o22a_1
XANTENNA__14260__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18325_ net599 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__inv_2
X_15537_ _01554_ _01555_ _01558_ _01469_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12749_ net501 _06620_ _06622_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__a21o_1
XANTENNA__11613__A2 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_332_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18256_ net644 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15468_ _08891_ _08892_ _01493_ _01494_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_170_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_301_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17207_ _02612_ net120 _02732_ net1698 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[485\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11589__A game.CPU.applesa.ab.check_walls.above.walls\[106\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14419_ game.CPU.applesa.ab.absxs.body_x\[111\] net874 net853 game.CPU.applesa.ab.absxs.body_y\[110\]
+ vssd1 vssd1 vccd1 vccd1 _08293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_331_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18187_ net608 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__inv_2
X_15399_ game.writer.updater.commands.count\[6\] game.writer.updater.commands.count\[5\]
+ _08888_ _01426_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__a31o_1
XFILLER_0_181_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_303_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19999__RESET_B net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12574__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17138_ _02405_ net72 net736 vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__o21a_1
Xhold604 game.writer.tracker.frame\[560\] vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09059__A game.CPU.applesa.ab.absxs.body_y\[52\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19917__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold615 game.writer.tracker.frame\[224\] vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 game.writer.tracker.frame\[21\] vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17501__A1 _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16451__Y _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold637 game.writer.tracker.frame\[392\] vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19928__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold648 game.writer.updater.commands.count\[13\] vssd1 vssd1 vccd1 vccd1 net2033
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11101__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17069_ net158 net82 vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__nand2_8
XANTENNA__12912__S net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold659 game.writer.tracker.frame\[5\] vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ net1155 _04188_ _04187_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_38_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13523__C1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09891_ _03613_ _03617_ _04064_ _04133_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkload19_A clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09506__B game.CPU.applesa.ab.absxs.body_y\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_191_Right_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_181_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17280__A3 _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13826__B1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10004__Y _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13743__S net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout184_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09522__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout351_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11852__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16240__A1 _06573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1093_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout449_A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14251__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16791__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_270_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09325_ net1105 _03266_ game.CPU.applesa.ab.absxs.body_y\[80\] net891 _03567_ vssd1
+ vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__o221a_1
XANTENNA__19447__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout616_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1358_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09256_ game.CPU.randy.counter1.count\[9\] vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__inv_2
XFILLER_0_334_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16074__B net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_322_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11499__A game.CPU.applesa.ab.check_walls.above.walls\[171\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09187_ game.CPU.applesa.ab.check_walls.above.walls\[104\] vssd1 vssd1 vccd1 vccd1
+ _03436_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16642__X _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1146_X net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19597__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13762__C1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16361__Y _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout985_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19669__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10040__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12107__B net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16846__A3 _02619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10591__A2 _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ _04283_ _04299_ _04307_ _04265_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__o211a_1
XANTENNA__16521__C _02373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13514__C1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_281_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11946__B net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11080_ game.CPU.applesa.ab.absxs.body_x\[43\] net544 net538 game.CPU.applesa.ab.absxs.body_y\[42\]
+ _04966_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__a221o_1
XFILLER_0_219_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10031_ net1134 _04237_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__and2_1
XANTENNA__09416__B game.CPU.applesa.ab.absxs.body_x\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15137__C game.CPU.applesa.ab.check_walls.above.walls\[165\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17008__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19902__Q game.writer.tracker.frame\[497\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13506__X _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13653__S net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14976__C net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14770_ game.CPU.randy.counter1.count\[6\] game.CPU.randy.counter1.count\[5\] game.CPU.randy.counter1.count\[8\]
+ game.CPU.randy.counter1.count\[7\] vssd1 vssd1 vccd1 vccd1 _08591_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11982_ game.CPU.applesa.ab.check_walls.above.walls\[181\] net388 vssd1 vssd1 vccd1
+ vccd1 _05869_ sky130_fd_sc_hd__xnor2_1
X_13721_ game.writer.tracker.frame\[198\] net843 net837 game.writer.tracker.frame\[197\]
+ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_205_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11681__B net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10933_ game.CPU.applesa.ab.absxs.body_y\[10\] net401 vssd1 vssd1 vccd1 vccd1 _04823_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_279_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ _02227_ _02400_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13045__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13652_ game.writer.tracker.frame\[33\] game.writer.tracker.frame\[35\] game.writer.tracker.frame\[36\]
+ game.writer.tracker.frame\[34\] net969 net1003 vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__mux4_1
X_10864_ _04749_ _04759_ _04761_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_292_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16782__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14992__B net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_143_Left_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_234_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11056__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12603_ game.CPU.applesa.ab.absxs.body_x\[93\] net375 vssd1 vssd1 vccd1 vccd1 _06480_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__13889__A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16371_ net134 _02259_ _02351_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__or3b_1
XFILLER_0_155_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13583_ _07455_ _07456_ net502 vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__mux2_1
X_10795_ game.CPU.applesa.ab.absxs.body_y\[42\] _04690_ _04728_ game.CPU.applesa.ab.absxs.body_y\[38\]
+ vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__a22o_1
XANTENNA__16265__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18110_ net632 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15322_ game.CPU.applesa.twomode.number\[1\] _08861_ net757 vssd1 vssd1 vccd1 vccd1
+ _08867_ sky130_fd_sc_hd__a21oi_1
XANTENNA__18814__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19090_ net1177 _00127_ _00761_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[135\]
+ sky130_fd_sc_hd__dfrtp_4
X_12534_ _06406_ _06408_ _06410_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__and3b_1
XFILLER_0_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18041_ net659 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_313_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15253_ game.CPU.kyle.L1.nextState\[4\] _08809_ net264 net2024 vssd1 vssd1 vccd1
+ vccd1 _01265_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12465_ game.CPU.applesa.ab.absxs.body_x\[15\] net530 vssd1 vssd1 vccd1 vccd1 _06342_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__12556__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_293_Right_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14204_ _03269_ net1075 net854 game.CPU.applesa.ab.absxs.body_y\[66\] _08075_ vssd1
+ vssd1 vccd1 vccd1 _08078_ sky130_fd_sc_hd__a221o_1
X_11416_ net775 _05304_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15184_ _04614_ _08752_ _08759_ game.CPU.bodymain1.main.score\[7\] vssd1 vssd1 vccd1
+ vccd1 _08760_ sky130_fd_sc_hd__o22a_1
XANTENNA__09421__B1 game.CPU.applesa.ab.absxs.body_x\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12396_ _06263_ _06265_ _06266_ _06267_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__or4_1
XANTENNA__12017__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11347_ game.CPU.applesa.ab.check_walls.above.walls\[139\] net760 vssd1 vssd1 vccd1
+ vccd1 _05236_ sky130_fd_sc_hd__xor2_2
XFILLER_0_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09972__A1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15609__A game.CPU.applesa.ab.absxs.body_y\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14135_ net887 game.CPU.applesa.ab.check_walls.above.walls\[40\] game.CPU.applesa.ab.check_walls.above.walls\[47\]
+ net857 vssd1 vssd1 vccd1 vccd1 _08009_ sky130_fd_sc_hd__a22o_1
XANTENNA__12732__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19992_ clknet_leaf_45_clk _01416_ net1299 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10582__A2 _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_152_Left_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11278_ _04974_ _04975_ _05166_ _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__or4b_1
X_14066_ net1058 game.CPU.applesa.ab.check_walls.above.walls\[2\] vssd1 vssd1 vccd1
+ vccd1 _07940_ sky130_fd_sc_hd__xnor2_1
X_18943_ net1176 _00082_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number_out\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11856__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_245_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09724__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13017_ game.writer.tracker.frame\[544\] game.writer.tracker.frame\[545\] net1021
+ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__mux2_1
X_10229_ game.CPU.applesa.ab.count_luck\[4\] game.CPU.applesa.ab.count_luck\[5\] _04421_
+ _04419_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__a31o_1
XANTENNA__09724__B2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18874_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[4\] _00569_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[4\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12033__A game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_342_Left_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17825_ game.writer.updater.commands.count\[3\] _03153_ vssd1 vssd1 vccd1 vccd1 _03157_
+ sky130_fd_sc_hd__or2_1
Xhold1 game.writer.control.button5.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_146_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17756_ _03112_ _03113_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14968_ net1272 _08744_ vssd1 vssd1 vccd1 vccd1 _08745_ sky130_fd_sc_hd__and2_1
XFILLER_0_221_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16707_ _02489_ net63 _02568_ net1841 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[149\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11591__B net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13919_ net1043 game.CPU.applesa.ab.check_walls.above.walls\[155\] vssd1 vssd1 vccd1
+ vccd1 _07793_ sky130_fd_sc_hd__or2_1
XANTENNA__15063__B net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17687_ _03062_ _03070_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_334_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14899_ _08674_ _08675_ vssd1 vssd1 vccd1 vccd1 _08676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_161_Left_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19426_ clknet_leaf_41_clk game.writer.tracker.next_frame\[21\] net1330 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_336_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13036__A1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16638_ net67 _02518_ _02537_ net1609 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[111\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16773__A2 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_256_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13799__A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_312_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19357_ clknet_leaf_70_clk game.CPU.applesa.twoapples.absxs.next_head\[2\] vssd1
+ vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.x_final\[2\] sky130_fd_sc_hd__dfxtp_1
X_16569_ net195 _02439_ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__nand2_2
X_09110_ net1434 vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__inv_2
X_18308_ net621 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_351_Left_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19288_ clknet_leaf_69_clk net403 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.y_final\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_304_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10935__B net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09041_ game.CPU.applesa.ab.absxs.body_x\[10\] vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__inv_2
XANTENNA__14407__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18239_ net650 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
XANTENNA__15733__B1 game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18390__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__A1_N net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13744__C1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_260_Right_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold401 game.CPU.randy.f1.c1.count\[14\] vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_276_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold412 game.writer.tracker.frame\[259\] vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_345_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold423 game.writer.tracker.frame\[395\] vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19762__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold434 game.writer.tracker.frame\[95\] vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09963__A1 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold445 game.writer.tracker.frame\[414\] vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 game.writer.tracker.frame\[149\] vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold467 game.writer.tracker.frame\[247\] vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__A2 net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold478 game.writer.tracker.frame\[433\] vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09517__A net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold489 game.writer.tracker.frame\[463\] vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ game.CPU.bodymain1.main.score\[7\] _04180_ vssd1 vssd1 vccd1 vccd1 _01393_
+ sky130_fd_sc_hd__xnor2_1
Xfanout903 net905 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_209_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 net915 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_4
XFILLER_0_96_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout925 net928 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13039__A net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout936 net937 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_2
XANTENNA__09715__A1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09715__B2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09874_ _04111_ _04114_ _04115_ _04116_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__or4_1
Xfanout947 net950 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__buf_4
Xfanout958 net959 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_4
Xfanout969 net972 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1106_A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11522__B2 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13981__B net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17253__A3 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_271_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout187_X net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout566_A _04460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16461__A1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12597__B net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16069__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_356_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout733_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1096_X net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16764__A2 _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16356__Y _02341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11006__B net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15701__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout900_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1263_X net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09308_ net1102 game.CPU.applesa.ab.absxs.body_x\[53\] vssd1 vssd1 vccd1 vccd1 _03551_
+ sky130_fd_sc_hd__xor2_1
X_10580_ _04174_ _04581_ _04655_ _04658_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__a31o_4
XANTENNA_clkbuf_leaf_7_clk_X clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14317__B net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09239_ net1 vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__inv_2
XANTENNA__17909__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18987__CLK net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13735__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12250_ game.CPU.applesa.ab.check_walls.above.walls\[119\] net424 vssd1 vssd1 vccd1
+ vccd1 _06136_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09403__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16532__B _02303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__A1 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ _03250_ net321 vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_309_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09954__A1 _03527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13750__A2 game.writer.tracker.frame\[144\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ _05868_ _05886_ _05950_ _06067_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.below.collision
+ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_151_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14333__A game.CPU.applesa.ab.absxs.body_x\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10564__A2 _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ game.CPU.applesa.ab.absxs.body_x\[69\] net322 vssd1 vssd1 vccd1 vccd1 _05022_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__09427__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15148__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11063_ game.CPU.applesa.ab.absxs.body_y\[24\] net533 vssd1 vssd1 vccd1 vccd1 _04953_
+ sky130_fd_sc_hd__nand2_1
X_15940_ game.CPU.applesa.ab.check_walls.above.walls\[43\] net458 vssd1 vssd1 vccd1
+ vccd1 _01952_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_275_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12710__B1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ net891 _04220_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__xnor2_2
XANTENNA__17244__A3 _02357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15871_ _03280_ net350 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_290_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16452__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19612__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17610_ _03021_ _03022_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__nor2_1
X_14822_ game.CPU.randy.counter1.count\[16\] _08626_ vssd1 vssd1 vccd1 vccd1 _08628_
+ sky130_fd_sc_hd__nand2_1
X_18590_ clknet_leaf_31_clk _01010_ _00327_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[59\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_188_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_240_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_230_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11277__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17541_ _03217_ _02772_ _02774_ _02967_ _03219_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__a32o_1
XANTENNA__13361__S1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14753_ _08575_ _08576_ net55 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__and3b_1
X_11965_ _05781_ _05852_ _05791_ _05809_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ game.writer.tracker.frame\[497\] game.writer.tracker.frame\[499\] game.writer.tracker.frame\[500\]
+ game.writer.tracker.frame\[498\] net975 net1014 vssd1 vssd1 vccd1 vccd1 _07578_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_230_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13018__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10916_ _04394_ _04472_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__or2_1
X_17472_ _02885_ _02899_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13018__B2 _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14215__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14684_ game.CPU.randy.counter1.count1\[9\] _08500_ _08504_ game.CPU.randy.counter1.count1\[8\]
+ _08522_ vssd1 vssd1 vccd1 vccd1 _08523_ sky130_fd_sc_hd__o221a_1
XANTENNA__16755__A2 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19762__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ net820 net312 vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__xnor2_1
X_19211_ net1167 _00023_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_possible\[2\]
+ sky130_fd_sc_hd__dfxtp_4
X_16423_ net195 _02347_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__nor2_8
X_13635_ game.writer.tracker.frame\[22\] net845 net838 game.writer.tracker.frame\[21\]
+ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__o22a_1
XANTENNA__13569__A2 game.writer.tracker.frame\[336\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10847_ _04747_ _04749_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_345_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19142_ net1184 _00184_ _00813_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[187\]
+ sky130_fd_sc_hd__dfrtp_4
X_16354_ _08028_ _02249_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__nand2_1
X_13566_ game.writer.tracker.frame\[365\] game.writer.tracker.frame\[367\] game.writer.tracker.frame\[368\]
+ game.writer.tracker.frame\[366\] net967 net997 vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__mux4_1
X_10778_ _04720_ game.CPU.applesa.ab.absxs.body_y\[59\] net327 vssd1 vssd1 vccd1 vccd1
+ _01010_ sky130_fd_sc_hd__mux2_1
XANTENNA__19079__Q game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_298_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14227__B net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15305_ game.CPU.applesa.twomode.counter _08849_ _08850_ _08851_ _08852_ vssd1 vssd1
+ vccd1 vccd1 _08853_ sky130_fd_sc_hd__a32o_1
XFILLER_0_109_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19073_ net1185 _00108_ _00744_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12517_ game.CPU.applesa.ab.absxs.body_y\[69\] net524 vssd1 vssd1 vccd1 vccd1 _06394_
+ sky130_fd_sc_hd__xnor2_1
X_16285_ game.writer.tracker.frame\[8\] net718 _02281_ _02287_ net135 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.next_frame\[8\] sky130_fd_sc_hd__a32o_1
X_13497_ _07061_ _07062_ net705 vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_297_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12529__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16133__A1_N game.CPU.applesa.ab.absxs.body_x\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13726__C1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_251_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18024_ net663 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15236_ _08797_ _08798_ _00019_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_340_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12448_ game.CPU.applesa.ab.absxs.body_x\[89\] net375 vssd1 vssd1 vccd1 vccd1 _06325_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_288_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18711__Q game.CPU.applesa.ab.absxs.body_x\[73\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15167_ net1226 net1253 game.CPU.walls.rand_wall.x_final\[3\] vssd1 vssd1 vccd1 vccd1
+ _00221_ sky130_fd_sc_hd__and3_1
XFILLER_0_288_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12379_ game.CPU.applesa.ab.absxs.body_y\[112\] net362 net369 _03323_ vssd1 vssd1
+ vccd1 vccd1 _06256_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12315__X _06201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19142__CLK net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14118_ net1043 _03472_ game.CPU.applesa.ab.check_walls.above.walls\[173\] net862
+ _07991_ vssd1 vssd1 vccd1 vccd1 _07992_ sky130_fd_sc_hd__a221o_1
XANTENNA__09337__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15058__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11586__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16140__B1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19975_ clknet_leaf_41_clk game.writer.tracker.next_frame\[570\] net1330 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[570\] sky130_fd_sc_hd__dfrtp_1
X_15098_ net1205 net1229 net794 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10490__B _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16691__A1 _02303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14049_ net959 game.CPU.applesa.ab.check_walls.above.walls\[197\] vssd1 vssd1 vccd1
+ vccd1 _07923_ sky130_fd_sc_hd__xor2_1
X_18926_ clknet_leaf_5_clk net1396 _00610_ vssd1 vssd1 vccd1 vccd1 game.CPU.right_button.eD1.Q1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_165_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_340_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17235__A3 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19292__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18857_ clknet_leaf_0_clk _01248_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19191__D net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15074__A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17808_ game.writer.updater.commands.cmd_num\[0\] _01436_ game.writer.updater.commands.cmd_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__or3b_1
X_09590_ net1094 _03388_ net827 net909 vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__o22a_1
X_18788_ clknet_leaf_9_clk _01203_ _00525_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_173_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14454__B1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17739_ _03101_ _03103_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__and2_1
XANTENNA__13352__S1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12210__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18385__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10011__A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16746__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14206__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09881__B1 _03774_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19409_ clknet_leaf_48_clk game.writer.tracker.next_frame\[4\] net1295 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[4\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15521__B net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10946__A game.CPU.applesa.ab.absxs.body_y\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout147_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_176_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_351_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_323_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10665__B _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout314_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17171__A2 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1056_A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10794__A2 _04690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ game.CPU.applesa.ab.absxs.body_x\[48\] vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__inv_2
XFILLER_0_331_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_248_Left_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11056__A1_N game.CPU.applesa.ab.absxs.body_y\[106\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold220 game.writer.tracker.frame\[203\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13732__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15249__A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout102_X net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold231 game.writer.tracker.frame\[487\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_198_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14153__A _08015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 game.writer.tracker.frame\[479\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_269_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1223_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold253 game.writer.tracker.frame\[154\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_269_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold264 game.writer.tracker.frame\[440\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold275 game.writer.tracker.frame\[145\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 game.writer.tracker.frame\[249\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout683_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout700 net701 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_4
Xhold297 game.writer.tracker.frame\[543\] vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout711 net712 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_4
XANTENNA__19635__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13992__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout722 net724 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_2
XANTENNA__16682__B2 _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09926_ _04148_ _04149_ net1109 vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a21o_1
Xfanout733 net738 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_2
XFILLER_0_284_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_187_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout744 net745 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1109_X net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20046_ game.CPU.randy.counter1.out vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
Xfanout766 net767 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09857_ net1094 game.CPU.applesa.ab.absxs.body_x\[46\] vssd1 vssd1 vccd1 vccd1 _04100_
+ sky130_fd_sc_hd__xnor2_1
Xfanout777 net778 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_304_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout788 game.CPU.applesa.ab.check_walls.above.walls\[159\] vssd1 vssd1 vccd1 vccd1
+ net788 sky130_fd_sc_hd__buf_2
XANTENNA_fanout471_X net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 game.CPU.applesa.ab.check_walls.above.walls\[116\] vssd1 vssd1 vccd1 vccd1
+ net799 sky130_fd_sc_hd__buf_2
XANTENNA_fanout569_X net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_257_Left_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09788_ _04021_ _04024_ _04025_ _04030_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__or4_1
XANTENNA__14445__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19785__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16985__A2 _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11259__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12120__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_233_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_202_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11750_ _03474_ net310 vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_68_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_276_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_218_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ game.CPU.applesa.ab.absxs.body_y\[77\] _04623_ _04624_ game.CPU.applesa.ab.absxs.body_y\[73\]
+ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__a22o_1
XFILLER_0_327_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ game.CPU.applesa.ab.check_walls.above.walls\[57\] net772 vssd1 vssd1 vccd1
+ vccd1 _05570_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14328__A game.CPU.applesa.ab.absxs.body_x\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_313_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13420_ _06993_ _07008_ net676 vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10632_ _03241_ net328 vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__nor2_1
XANTENNA__15150__C game.CPU.applesa.ab.check_walls.above.walls\[178\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_342_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12854__S0 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13351_ net226 _07223_ net283 vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__a21o_1
X_10563_ net1080 _04653_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_153_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17162__A2 _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_279_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_266_Left_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19165__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12302_ _05903_ _06187_ _05905_ _05904_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__or4bb_1
X_16070_ game.CPU.applesa.ab.absxs.body_x\[86\] net346 vssd1 vssd1 vccd1 vccd1 _02082_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13282_ _07153_ _07154_ net683 vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__mux2_1
X_10494_ _03197_ net1120 vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__nor2_1
XFILLER_0_295_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15021_ net1222 net1250 game.CPU.applesa.ab.check_walls.above.walls\[49\] vssd1 vssd1
+ vccd1 vccd1 _00240_ sky130_fd_sc_hd__and3_1
XANTENNA__13723__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_267_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15159__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12233_ net814 net420 vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_287_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11734__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10537__A2 _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ _05523_ _05526_ _06050_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__or3_1
XANTENNA__09157__A game.CPU.applesa.ab.check_walls.above.walls\[49\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16122__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_229_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11115_ _04999_ _05001_ _05002_ _05003_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__or4_1
X_16972_ _02445_ _02638_ net730 vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__o21a_1
X_19760_ clknet_leaf_26_clk game.writer.tracker.next_frame\[355\] net1313 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[355\] sky130_fd_sc_hd__dfrtp_1
X_12095_ _05981_ _05980_ _05979_ _05978_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__and4b_1
XANTENNA__13487__A1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17805__C _06573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18711_ clknet_leaf_60_clk _01128_ _00448_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[73\]
+ sky130_fd_sc_hd__dfrtp_4
X_15923_ game.CPU.applesa.ab.check_walls.above.walls\[130\] net346 vssd1 vssd1 vccd1
+ vccd1 _01935_ sky130_fd_sc_hd__nand2_1
X_11046_ _03266_ net326 vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__xnor2_2
X_19691_ clknet_leaf_25_clk game.writer.tracker.next_frame\[286\] net1320 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[286\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17217__A3 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_275_Left_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16425__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18642_ clknet_leaf_53_clk _01059_ _00379_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[44\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_290_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15854_ _03262_ net270 vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_274_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14436__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14805_ _08616_ _08617_ vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18573_ clknet_leaf_62_clk _00993_ _00310_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_15785_ game.CPU.applesa.ab.absxs.body_y\[74\] net335 vssd1 vssd1 vccd1 vccd1 _01797_
+ sky130_fd_sc_hd__nand2_1
X_12997_ game.writer.tracker.frame\[518\] game.writer.tracker.frame\[519\] net1008
+ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16718__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17524_ _02841_ _02950_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__nand2_1
X_14736_ _03502_ _08563_ vssd1 vssd1 vccd1 vccd1 _08565_ sky130_fd_sc_hd__nor2_1
XANTENNA__16189__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ net748 _05302_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__nand2_1
XANTENNA__16728__A2 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_290_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11670__B1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17455_ _03197_ _02786_ _02787_ _02792_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__o22a_1
XFILLER_0_357_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15936__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14667_ game.CPU.randy.counter1.count1\[6\] _04348_ net266 vssd1 vssd1 vccd1 vccd1
+ _08506_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_253_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14238__A game.CPU.applesa.ab.absxs.body_x\[114\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11879_ game.CPU.applesa.ab.check_walls.above.walls\[141\] net305 net299 net791 vssd1
+ vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a22oi_1
X_16406_ _02262_ _02279_ _02333_ _01516_ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__a22oi_4
X_13618_ game.writer.tracker.frame\[281\] game.writer.tracker.frame\[283\] game.writer.tracker.frame\[284\]
+ game.writer.tracker.frame\[282\] net975 net1017 vssd1 vssd1 vccd1 vccd1 _07492_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_223_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13411__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19508__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17386_ game.CPU.kyle.L1.nextState\[5\] game.CPU.kyle.L1.nextState\[4\] vssd1 vssd1
+ vccd1 vccd1 _02816_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_284_Left_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14598_ game.CPU.clock1.counter\[3\] _08455_ _08456_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[3\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__16724__Y _02577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19125_ net1183 _00166_ _00796_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[170\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_333_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16337_ net136 _02278_ _02327_ _02324_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[20\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13549_ _07421_ _07422_ net478 vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__mux2_1
XANTENNA__16453__A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10776__A2 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19056_ net1191 _00090_ _00727_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[101\]
+ sky130_fd_sc_hd__dfrtp_1
X_16268_ net132 _02272_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__nand2_8
XTAP_TAPCELL_ROW_329_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16900__A2 _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18007_ net616 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__inv_2
XANTENNA__19658__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15219_ game.CPU.applesa.normal1.number\[0\] _08780_ vssd1 vssd1 vccd1 vccd1 _08785_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09918__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14911__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16199_ game.CPU.applesa.ab.absxs.body_x\[57\] net473 net462 game.CPU.applesa.ab.absxs.body_x\[59\]
+ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10528__A2 _04609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11725__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09067__A game.CPU.applesa.ab.absxs.body_y\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17310__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16664__B2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19958_ clknet_leaf_44_clk game.writer.tracker.next_frame\[553\] net1304 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[553\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10006__A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_293_Left_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_206_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18682__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12699__Y _06573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ net1139 game.CPU.applesa.ab.absxs.body_y\[22\] vssd1 vssd1 vccd1 vccd1 _03954_
+ sky130_fd_sc_hd__xor2_1
X_18909_ clknet_leaf_4_clk _01276_ _00593_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_19889_ clknet_leaf_27_clk game.writer.tracker.next_frame\[484\] net1309 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[484\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16416__A1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09642_ net1154 game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1 vccd1
+ vccd1 _03885_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16967__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10700__A2 _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09573_ net1088 game.CPU.applesa.ab.check_walls.above.walls\[43\] vssd1 vssd1 vccd1
+ vccd1 _03816_ sky130_fd_sc_hd__xor2_1
XFILLER_0_210_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_353_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13650__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10464__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_309_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout431_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1173_A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout529_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_351_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17144__A2 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1059_X net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__A2 _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13166__A0 _07032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_249_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16082__B net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout898_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09007_ game.CPU.applesa.ab.absxs.body_x\[112\] vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_189_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_276_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_249_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11716__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_306_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__A2 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16655__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13469__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_284_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout530 net532 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_4
Xfanout541 _04816_ vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__buf_4
Xfanout552 net555 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_2
X_09909_ net1092 _04147_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__xnor2_1
Xfanout563 net564 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout574 net575 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_232_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout585 net587 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_2
X_12920_ _06783_ _06788_ _06792_ _06793_ net247 vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__o221a_1
XFILLER_0_232_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout596 net598 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__buf_4
X_20029_ net1276 vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
XANTENNA__15145__C game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16958__A2 _02415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_224_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17080__A1 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12851_ game.writer.tracker.frame\[268\] game.writer.tracker.frame\[269\] net996
+ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16422__A4 _02387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16538__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15630__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11802_ net816 net313 vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14984__C game.CPU.applesa.ab.check_walls.above.walls\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15570_ net1416 net1419 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__xnor2_1
X_12782_ game.writer.tracker.frame\[90\] game.writer.tracker.frame\[91\] net1019 vssd1
+ vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__mux2_1
XANTENNA__12444__A2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14521_ _08040_ _08369_ _08393_ vssd1 vssd1 vccd1 vccd1 _08395_ sky130_fd_sc_hd__and3b_1
X_11733_ net570 _05476_ _05481_ _05482_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__o211a_1
XANTENNA__14058__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17240_ net157 _02432_ net72 net729 vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__o31a_1
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14452_ game.CPU.applesa.ab.absxs.body_x\[12\] net1074 vssd1 vssd1 vccd1 vccd1 _08326_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11664_ game.CPU.applesa.ab.check_walls.above.walls\[120\] net773 vssd1 vssd1 vccd1
+ vccd1 _05553_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_315_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13403_ _07275_ _07276_ net484 vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__mux2_1
XANTENNA__18555__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17171_ net147 _02467_ net73 _02723_ net1470 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[458\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__11404__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10615_ game.CPU.applesa.ab.absxs.body_x\[74\] _04675_ _04676_ game.CPU.applesa.ab.absxs.body_x\[70\]
+ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_289_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13944__A2 game.CPU.applesa.ab.check_walls.above.walls\[68\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14383_ _03266_ net1069 net947 _03329_ _08252_ vssd1 vssd1 vccd1 vccd1 _08257_ sky130_fd_sc_hd__o221a_1
XANTENNA__19800__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17135__A2 _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11595_ game.CPU.applesa.ab.check_walls.above.walls\[109\] net315 vssd1 vssd1 vccd1
+ vccd1 _05484_ sky130_fd_sc_hd__nand2_1
X_16122_ game.CPU.applesa.ab.absxs.body_x\[54\] net467 net441 game.CPU.applesa.ab.absxs.body_y\[54\]
+ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13334_ net219 _07204_ _07207_ net282 vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__a211o_1
X_10546_ net848 _04644_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__or2_4
XANTENNA__15697__A2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16894__A1 _02464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16053_ _03227_ net349 net335 _03293_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__a22o_1
X_13265_ game.writer.tracker.frame\[486\] game.writer.tracker.frame\[487\] net999
+ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__mux2_1
XANTENNA__10525__S _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10477_ _03264_ _04601_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__nor2_1
X_15004_ net1221 net1249 game.CPU.applesa.ab.check_walls.above.walls\[32\] vssd1 vssd1
+ vccd1 vccd1 _00222_ sky130_fd_sc_hd__and3_1
XFILLER_0_283_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12216_ game.CPU.applesa.ab.check_walls.above.walls\[5\] net549 vssd1 vssd1 vccd1
+ vccd1 _06102_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19950__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13196_ _07066_ _07067_ _07069_ _07068_ net497 net689 vssd1 vssd1 vccd1 vccd1 _07070_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_283_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_282_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12380__A1 game.CPU.applesa.ab.absxs.body_y\[113\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19812_ clknet_leaf_37_clk game.writer.tracker.next_frame\[407\] net1351 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[407\] sky130_fd_sc_hd__dfrtp_1
X_12147_ _06031_ _06032_ _06033_ _06026_ _06020_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__o311a_1
XFILLER_0_263_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_263_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09615__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19743_ clknet_leaf_25_clk game.writer.tracker.next_frame\[338\] net1341 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[338\] sky130_fd_sc_hd__dfrtp_1
X_16955_ _02410_ net94 _02657_ net1811 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[308\]
+ sky130_fd_sc_hd__a22o_1
X_12078_ net808 net294 vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__nand2_1
XANTENNA__12132__A1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12132__B2 game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15906_ _03339_ net337 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__xnor2_1
X_11029_ _03269_ net415 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__nand2_1
X_16886_ net1878 _02631_ net97 _02454_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[260\]
+ sky130_fd_sc_hd__a22o_1
X_19674_ clknet_leaf_32_clk game.writer.tracker.next_frame\[269\] net1285 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[269\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15055__C game.CPU.applesa.ab.check_walls.above.walls\[83\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16949__A2 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13880__A1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14409__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13880__B2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17071__A1 _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__X _04145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15837_ game.CPU.applesa.ab.check_walls.above.walls\[18\] net348 vssd1 vssd1 vccd1
+ vccd1 _01849_ sky130_fd_sc_hd__nand2_1
X_18625_ clknet_leaf_11_clk _01042_ _00362_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[107\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16448__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13571__S net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15768_ _03288_ net272 net341 _03355_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__a22o_1
X_18556_ clknet_leaf_1_clk _00012_ net429 vssd1 vssd1 vccd1 vccd1 game.CPU.speed1.Qa\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_59_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19330__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17507_ net1264 _02837_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__nor2_1
X_14719_ game.CPU.randy.counter1.count1\[5\] _08551_ vssd1 vssd1 vccd1 vccd1 _08554_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18487_ net631 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15699_ _01703_ _01706_ _01707_ _01708_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__or4_1
XFILLER_0_318_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_318_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17438_ _02781_ _02815_ _02865_ _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a211o_1
XFILLER_0_129_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_318_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_32_clk_X clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 _04118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_26 _07032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16454__Y _02412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 game.writer.tracker.frame\[113\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_48 game.writer.tracker.frame\[305\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11104__B net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19480__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17369_ _02798_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__inv_2
XANTENNA__12915__S net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14255__X _08129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17126__A2 _02382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10749__A2 _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19108_ net1180 _00147_ _00779_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[153\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10943__B net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload49_A clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_47_clk_X clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19039_ net1189 _00270_ _00710_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_286_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16885__B2 _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_212_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16470__X _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13699__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09509__B game.CPU.applesa.ab.absxs.body_y\[50\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12216__A game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14360__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16637__A1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_329_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15663__A2_N game.CPU.applesa.ab.check_walls.above.walls\[55\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout381_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12123__A1 game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout479_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12123__B2 game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_301_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_254_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_345_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17062__A1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09625_ _03861_ _03863_ _03866_ _03867_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__or4_2
XANTENNA__11882__B1 _05769_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1290_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout646_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09556_ net917 game.CPU.applesa.ab.absxs.body_x\[61\] game.CPU.applesa.ab.absxs.body_x\[60\]
+ net913 vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__a22o_1
XFILLER_0_328_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16077__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_273_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09487_ net1126 net781 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19823__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16573__B1 _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_352_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_336_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_230_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1343_X net1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_312_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17117__A2 _02693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_199_Left_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10400_ _04547_ _04549_ _04341_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__o21ai_1
X_11380_ net775 _05268_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19973__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14325__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10331_ game.CPU.randy.f1.a1.count\[7\] _04490_ game.CPU.randy.f1.a1.count\[8\] vssd1
+ vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a21o_1
XANTENNA__17917__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09419__B game.CPU.applesa.ab.absxs.body_y\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_249_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13050_ game.writer.tracker.frame\[256\] game.writer.tracker.frame\[257\] net1032
+ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__mux2_2
XFILLER_0_265_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10262_ _04452_ _04454_ _04449_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__a21o_1
XFILLER_0_249_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_284_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16540__B _02311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19203__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13656__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12001_ game.CPU.applesa.ab.check_walls.above.walls\[164\] net552 vssd1 vssd1 vccd1
+ vccd1 _05888_ sky130_fd_sc_hd__nand2_1
XANTENNA__13509__X _07383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_226_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10193_ _04384_ _04385_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout82_X net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1303 net1305 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__clkbuf_4
Xfanout1314 net1360 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__clkbuf_2
Xfanout1325 net1334 vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09435__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1336 net1337 vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__buf_2
XANTENNA__15156__B net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1347 net1348 vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_148_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1358 net1359 vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__clkbuf_2
Xfanout360 net362 vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__buf_4
Xfanout371 net374 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_4
XFILLER_0_260_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16740_ _02375_ net61 _02582_ net1673 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[168\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout382 net385 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_4
XFILLER_0_255_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13952_ _07824_ _07825_ vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__nand2_1
Xfanout393 net394 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_260_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19353__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17053__A1 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12903_ game.writer.tracker.frame\[22\] game.writer.tracker.frame\[23\] net1024 vssd1
+ vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16671_ net2007 _02550_ _02553_ net127 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[128\]
+ sky130_fd_sc_hd__a22o_1
X_13883_ net1055 game.CPU.applesa.ab.check_walls.above.walls\[98\] vssd1 vssd1 vccd1
+ vccd1 _07757_ sky130_fd_sc_hd__xor2_1
XANTENNA__16268__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16800__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15622_ game.CPU.applesa.ab.absxs.body_y\[71\] net435 vssd1 vssd1 vccd1 vccd1 _01634_
+ sky130_fd_sc_hd__xnor2_1
X_18410_ net602 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__inv_2
X_12834_ _06704_ _06705_ _06707_ _06706_ net490 net683 vssd1 vssd1 vccd1 vccd1 _06708_
+ sky130_fd_sc_hd__mux4_1
X_19390_ clknet_leaf_8_clk _01396_ _00970_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.snake_head_x\[2\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_0_347_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_295_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09170__A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18341_ net595 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15553_ _01475_ _01572_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_29_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _06632_ _06633_ _06635_ _06637_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__or4_2
XANTENNA__09294__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_237_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09294__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14504_ game.CPU.apple_location\[7\] net856 net947 _03208_ vssd1 vssd1 vccd1 vccd1
+ _08378_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18272_ net664 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
X_11716_ net569 _04776_ _05603_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__o21ai_1
X_15484_ net888 _01505_ _01507_ net871 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__o22a_1
X_12696_ net1076 net955 vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__or2_2
XFILLER_0_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16715__B _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13378__B1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17223_ _02538_ net75 _02736_ game.writer.tracker.frame\[497\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[497\] sky130_fd_sc_hd__a22o_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14435_ game.CPU.applesa.ab.absxs.body_x\[27\] net876 net863 game.CPU.applesa.ab.absxs.body_y\[25\]
+ vssd1 vssd1 vccd1 vccd1 _08309_ sky130_fd_sc_hd__a22o_1
XANTENNA__13917__A2 game.CPU.applesa.ab.check_walls.above.walls\[157\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11647_ net777 _05535_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17108__A2 _02351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11928__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17154_ _02432_ _02693_ net736 vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__o21a_1
XANTENNA__16434__C _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14366_ _08239_ _08231_ _08234_ vssd1 vssd1 vccd1 vccd1 _08240_ sky130_fd_sc_hd__or3b_1
X_11578_ net563 _05459_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__nand2_1
XANTENNA__16867__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16105_ _01841_ _01842_ _02114_ _02115_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a22o_1
X_13317_ net490 _06729_ _07190_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10600__A1 game.CPU.applesa.ab.absxs.body_x\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17085_ _02309_ net57 _02697_ net1908 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[398\]
+ sky130_fd_sc_hd__a22o_1
X_10529_ game.CPU.applesa.ab.absxs.body_x\[53\] _04609_ _04637_ net1269 vssd1 vssd1
+ vccd1 vccd1 _01176_ sky130_fd_sc_hd__a22o_1
X_14297_ game.CPU.applesa.ab.absxs.body_x\[55\] net874 net964 _03307_ _08170_ vssd1
+ vssd1 vccd1 vccd1 _08171_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_326_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16036_ game.CPU.applesa.ab.absxs.body_y\[47\] net434 vssd1 vssd1 vccd1 vccd1 _02048_
+ sky130_fd_sc_hd__and2_1
X_13248_ game.writer.tracker.frame\[472\] game.writer.tracker.frame\[473\] net1016
+ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__mux2_1
XANTENNA__14342__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_256_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_248_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16619__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11875__A game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ game.writer.tracker.frame\[416\] game.writer.tracker.frame\[417\] net1037
+ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_296_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17292__A1 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17987_ net634 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__inv_2
XANTENNA__12105__B2 game.CPU.applesa.ab.check_walls.above.walls\[119\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19726_ clknet_leaf_22_clk game.writer.tracker.next_frame\[321\] net1342 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[321\] sky130_fd_sc_hd__dfrtp_1
X_16938_ _02375_ net92 _02652_ net1577 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[296\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13853__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17044__A1 _02404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19657_ clknet_leaf_22_clk game.writer.tracker.next_frame\[252\] net1347 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[252\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_315_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10667__B2 game.CPU.applesa.ab.absxs.body_x\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16869_ net153 _02424_ net107 _02628_ net1748 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[251\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__18720__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_337_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09410_ net891 net793 game.CPU.applesa.ab.check_walls.above.walls\[135\] net906 _03648_
+ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__a221o_1
XANTENNA__15082__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18608_ clknet_leaf_70_clk _01025_ _00345_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[90\]
+ sky130_fd_sc_hd__dfrtp_4
X_19588_ clknet_leaf_36_clk game.writer.tracker.next_frame\[183\] net1351 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[183\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13605__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_259_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09341_ net898 game.CPU.applesa.ab.absxs.body_y\[89\] game.CPU.applesa.ab.absxs.body_y\[88\]
+ net892 _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a221o_1
X_18539_ net612 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_331_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09272_ game.CPU.clock1.counter\[17\] vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18870__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19996__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14030__A1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14030__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11919__A1 game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout227_A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16344__C net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11769__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16858__A1 _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_348_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_259_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1136_A net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15530__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_302_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_247_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19725__Q game.writer.tracker.frame\[320\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13541__A0 game.writer.tracker.frame\[113\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16360__B _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout596_A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13476__S net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11785__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19376__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17283__A1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09760__A2 game.CPU.applesa.ab.check_walls.above.walls\[26\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout763_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ game.CPU.applesa.ab.absxs.body_x\[77\] vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12647__A2 game.CPU.applesa.twoapples.absxs.next_head\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16359__Y _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17035__A1 _02299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11009__B net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15704__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10658__B2 game.CPU.applesa.ab.absxs.body_x\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_230_Left_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout930_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1293_X net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_221_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16389__A3 _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09608_ net1111 game.CPU.applesa.ab.absxs.body_x\[116\] vssd1 vssd1 vccd1 vccd1 _03851_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_329_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10880_ game.CPU.applesa.ab.apple_possible\[7\] _04780_ vssd1 vssd1 vccd1 vccd1 _04782_
+ sky130_fd_sc_hd__xor2_4
XFILLER_0_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09539_ net1108 _03421_ game.CPU.applesa.ab.check_walls.above.walls\[76\] net892
+ _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_305_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_274_Right_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_241_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12550_ game.CPU.applesa.ab.absxs.body_y\[22\] net518 vssd1 vssd1 vccd1 vccd1 _06427_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ net564 _05388_ _05387_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_324_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12481_ game.CPU.applesa.ab.absxs.body_y\[29\] net523 net359 game.CPU.applesa.ab.absxs.body_y\[28\]
+ _06357_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12170__A1_N net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16561__A3 _02322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13240__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14220_ _03344_ net986 net952 _03343_ _08093_ vssd1 vssd1 vccd1 vccd1 _08094_ sky130_fd_sc_hd__a221o_1
XFILLER_0_321_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11432_ game.CPU.applesa.ab.check_walls.above.walls\[26\] net768 vssd1 vssd1 vccd1
+ vccd1 _05321_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_163_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_340_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11679__B game.CPU.applesa.ab.apple_possible\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14055__B net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16849__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_232_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11386__A2 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13780__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151_ net942 net951 net840 _07766_ _07812_ vssd1 vssd1 vccd1 vccd1 _08025_ sky130_fd_sc_hd__o311a_2
X_11363_ net824 net252 net317 net823 vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ net212 _06942_ _06975_ net283 vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__a211o_1
XFILLER_0_277_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19719__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10314_ _04487_ _04496_ net739 vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__a21o_1
X_14082_ net1072 _03427_ net807 net869 _07954_ vssd1 vssd1 vccd1 vccd1 _07956_ sky130_fd_sc_hd__o221a_1
X_11294_ _04910_ _04911_ _04912_ _04917_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__or4_1
XANTENNA__13532__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13386__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13033_ net484 _06904_ _06906_ net281 vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__a211o_1
XFILLER_0_265_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17910_ net662 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__inv_2
XFILLER_0_292_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_266_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10245_ _04418_ _04437_ _04416_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__a21o_1
XANTENNA__14071__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18890_ clknet_leaf_2_clk _01262_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1100 net1101 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__buf_4
XANTENNA__17274__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1111 net1112 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__buf_4
XANTENNA__09165__A game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17841_ game.writer.updater.commands.count\[8\] _01493_ _03158_ vssd1 vssd1 vccd1
+ vccd1 _03168_ sky130_fd_sc_hd__nand3_1
XANTENNA__09751__A2 game.CPU.applesa.ab.check_walls.above.walls\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ net1168 game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1 vccd1 vccd1 _04369_
+ sky130_fd_sc_hd__nand2_2
Xfanout1122 net1123 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__buf_1
XFILLER_0_206_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1133 game.CPU.applesa.ab.snake_head_y\[3\] vssd1 vssd1 vccd1 vccd1 net1133
+ sky130_fd_sc_hd__buf_4
XFILLER_0_280_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1144 net1152 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__buf_4
XANTENNA__12303__B net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18743__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19869__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1155 net1157 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_8
Xfanout1166 game.CPU.applesa.ab.logic_enable vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__buf_2
X_17772_ game.CPU.applesa.twoapples.count_luck\[7\] game.CPU.applesa.twoapples.count_luck\[6\]
+ _03121_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__nand3_1
Xfanout1177 net1178 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__buf_2
X_14984_ net1224 net1251 game.CPU.applesa.ab.check_walls.above.walls\[12\] vssd1 vssd1
+ vccd1 vccd1 _00200_ sky130_fd_sc_hd__and3_1
Xfanout190 net191 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__buf_4
Xfanout1188 net1189 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17026__A1 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16269__Y _02275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1199 net1201 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__clkbuf_2
X_19511_ clknet_leaf_14_clk game.writer.tracker.next_frame\[106\] net1283 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[106\] sky130_fd_sc_hd__dfrtp_1
X_16723_ net160 _02348_ net106 _02575_ net1715 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[157\]
+ sky130_fd_sc_hd__a32o_1
X_13935_ net951 net822 vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__xor2_1
XANTENNA__15614__B net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17577__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload5_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16654_ net152 _02419_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__nand2_1
X_19442_ clknet_leaf_47_clk game.writer.tracker.next_frame\[37\] net1299 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[37\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_282_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13866_ net225 _07710_ _07720_ _07739_ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_18_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15588__B2 game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15605_ net799 net449 net438 net797 _01616_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__a221o_1
X_12817_ game.writer.tracker.frame\[324\] game.writer.tracker.frame\[325\] net1030
+ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__mux2_1
X_16585_ net1780 _02500_ _02503_ net126 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[92\]
+ sky130_fd_sc_hd__a22o_1
X_19373_ clknet_leaf_70_clk _01379_ _00954_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location2\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_13797_ game.writer.tracker.frame\[387\] net710 net837 game.writer.tracker.frame\[385\]
+ vssd1 vssd1 vccd1 vccd1 _07671_ sky130_fd_sc_hd__o22a_1
XANTENNA__17329__A2 _02435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14260__A1 net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_241_Right_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15536_ _01544_ _01547_ _01556_ _01557_ _01553_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__o221a_1
X_18324_ net599 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__inv_2
X_12748_ net477 _06621_ net678 vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16445__B net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19249__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_343_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18255_ net645 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
XANTENNA__10821__A1 game.CPU.applesa.ab.absxs.body_y\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_154_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_332_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15467_ game.writer.updater.commands.count\[16\] game.writer.updater.commands.count\[9\]
+ game.writer.updater.commands.count\[8\] game.writer.updater.commands.count\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__or4b_1
X_12679_ _06551_ _06552_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14246__A game.CPU.applesa.ab.absxs.body_x\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17206_ _02611_ net120 _02732_ net1711 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[484\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_170_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14418_ game.CPU.applesa.ab.absxs.body_x\[108\] net1074 vssd1 vssd1 vccd1 vccd1 _08292_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11589__B net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18186_ net608 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__inv_2
XANTENNA__13220__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15398_ game.writer.updater.commands.count\[12\] game.writer.updater.commands.count\[9\]
+ game.writer.updater.commands.count\[8\] game.writer.updater.commands.count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__or4_1
XFILLER_0_114_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12574__A1 game.CPU.applesa.ab.absxs.body_y\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17137_ _02404_ net60 _02713_ net1542 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[434\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13771__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12574__B2 game.CPU.applesa.ab.absxs.body_y\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14349_ game.CPU.applesa.ab.absxs.body_x\[35\] net1045 vssd1 vssd1 vccd1 vccd1 _08223_
+ sky130_fd_sc_hd__xnor2_1
Xhold605 game.CPU.randy.f1.a1.count\[1\] vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 game.writer.tracker.frame\[340\] vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold627 game.writer.tracker.frame\[388\] vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19399__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold638 game.CPU.randy.f1.c1.count\[11\] vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 game.writer.tracker.frame\[448\] vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
X_17068_ net155 net72 vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__nor2_2
Xmax_cap357 _08416_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_4
XFILLER_0_311_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13296__S net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19194__D net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15077__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16019_ _03246_ net273 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_228_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09890_ _03623_ _03626_ _03566_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__o21a_1
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17265__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_271_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12213__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18388__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_264_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10014__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13287__C1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19709_ clknet_leaf_32_clk game.writer.tracker.next_frame\[304\] net1286 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[304\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09803__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11962__A1_N game.CPU.applesa.ab.check_walls.above.walls\[68\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_A _06639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16339__C _02328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09522__B game.CPU.applesa.ab.check_walls.above.walls\[123\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_338_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_338_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11490__D _05217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13685__S0 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16636__A net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout344_A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09324_ net902 game.CPU.applesa.ab.absxs.body_y\[82\] game.CPU.applesa.ab.absxs.body_y\[81\]
+ net897 vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_105_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_270_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_306_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_192_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09255_ game.CPU.randy.counter1.count\[10\] vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__inv_2
XANTENNA__18624__Q game.CPU.applesa.ab.absxs.body_y\[106\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout511_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13437__S0 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14156__A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14003__B2 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18616__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_322_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11499__B net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12014__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13211__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09186_ net802 vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__inv_2
XFILLER_0_321_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15539__X net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13995__A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16371__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1041_X net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09430__B2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1139_X net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16700__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18766__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout978_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_281_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1306_X net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17256__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ net1134 _04237_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__nor2_1
XFILLER_0_262_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_234_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18298__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_343_Right_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17008__A1 _02494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11981_ _05859_ _05862_ _05867_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__or3b_1
XFILLER_0_98_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13720_ game.writer.tracker.frame\[199\] net710 net673 game.writer.tracker.frame\[200\]
+ vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__o22a_1
XFILLER_0_242_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10932_ game.CPU.applesa.ab.absxs.body_y\[10\] net401 vssd1 vssd1 vccd1 vccd1 _04822_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_205_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15153__C game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_279_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10578__B net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13651_ game.writer.tracker.frame\[37\] game.writer.tracker.frame\[39\] game.writer.tracker.frame\[40\]
+ game.writer.tracker.frame\[38\] net970 net1003 vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__mux4_1
X_10863_ _04761_ _04762_ _04765_ _04740_ _04739_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_292_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16546__A net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15450__A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12602_ _06471_ _06472_ _06478_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__or3_1
XANTENNA__14992__C game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16370_ net197 _02350_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_26_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13582_ game.writer.tracker.frame\[373\] game.writer.tracker.frame\[375\] game.writer.tracker.frame\[376\]
+ game.writer.tracker.frame\[374\] net976 net1012 vssd1 vssd1 vccd1 vccd1 _07456_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_234_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ game.CPU.applesa.ab.absxs.body_y\[43\] _04690_ _04728_ game.CPU.applesa.ab.absxs.body_y\[39\]
+ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__a22o_1
XANTENNA__16265__B net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15321_ game.CPU.applesa.twomode.number\[1\] _08861_ vssd1 vssd1 vccd1 vccd1 _08866_
+ sky130_fd_sc_hd__or2_1
XANTENNA__19279__D game.CPU.applesa.ab.absxs.collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_183_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12533_ game.CPU.applesa.ab.absxs.body_x\[99\] net529 net518 game.CPU.applesa.ab.absxs.body_y\[98\]
+ _06409_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__o221a_1
XANTENNA__10803__A1 game.CPU.applesa.ab.absxs.body_y\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_81_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10803__B2 game.CPU.applesa.ab.absxs.body_y\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17192__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14066__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18040_ net613 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__inv_2
XANTENNA__12005__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15252_ _08812_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19541__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12464_ game.CPU.applesa.ab.absxs.body_x\[12\] net382 vssd1 vssd1 vccd1 vccd1 _06341_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14203_ game.CPU.applesa.ab.absxs.body_y\[64\] net870 net956 _03334_ vssd1 vssd1
+ vccd1 vccd1 _08077_ sky130_fd_sc_hd__a22o_1
XFILLER_0_297_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11415_ game.CPU.applesa.ab.check_walls.above.walls\[113\] net770 vssd1 vssd1 vccd1
+ vccd1 _05304_ sky130_fd_sc_hd__xor2_1
XANTENNA__11202__B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15183_ net1115 game.CPU.bodymain1.main.score\[4\] net1114 vssd1 vssd1 vccd1 vccd1
+ _08759_ sky130_fd_sc_hd__o21a_1
XANTENNA__09421__A1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12395_ _03280_ game.CPU.applesa.twoapples.absxs.next_head\[1\] game.CPU.applesa.twoapples.absxs.next_head\[6\]
+ _03349_ _06270_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__a221o_1
XFILLER_0_340_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09421__B2 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14134_ _08004_ _08005_ _08006_ _08007_ vssd1 vssd1 vccd1 vccd1 _08008_ sky130_fd_sc_hd__or4_1
X_11346_ game.CPU.applesa.ab.check_walls.above.walls\[138\] net765 vssd1 vssd1 vccd1
+ vccd1 _05235_ sky130_fd_sc_hd__xor2_2
XANTENNA__09972__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19991_ clknet_leaf_45_clk _01415_ net1304 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__15609__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14513__B net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19691__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14065_ net1068 game.CPU.applesa.ab.check_walls.above.walls\[1\] vssd1 vssd1 vccd1
+ vccd1 _07939_ sky130_fd_sc_hd__xnor2_1
X_18942_ net1176 _00081_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number_out\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11277_ game.CPU.applesa.ab.absxs.body_x\[61\] net412 net409 game.CPU.applesa.ab.absxs.body_x\[62\]
+ _04980_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_245_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13016_ game.writer.tracker.frame\[536\] game.writer.tracker.frame\[537\] net1022
+ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__mux2_1
XANTENNA__17247__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ game.CPU.applesa.ab.count_luck\[3\] _04420_ vssd1 vssd1 vccd1 vccd1 _04421_
+ sky130_fd_sc_hd__or2_1
X_18873_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[3\] _00568_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[3\] sky130_fd_sc_hd__dfrtp_1
X_17824_ game.writer.updater.commands.count\[3\] _03153_ vssd1 vssd1 vccd1 vccd1 _03156_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_310_Right_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2 game.CPU.down_button.eD1.D vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ _04343_ _04344_ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__or3_1
XANTENNA__18001__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17755_ game.CPU.applesa.twoapples.count_luck\[1\] game.CPU.applesa.twoapples.count_luck\[0\]
+ _03107_ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__and3_1
X_14967_ _08723_ _08740_ _08743_ _08733_ vssd1 vssd1 vccd1 vccd1 _08744_ sky130_fd_sc_hd__a31o_1
XFILLER_0_233_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16706_ _02327_ net63 _02568_ net1727 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[148\]
+ sky130_fd_sc_hd__a22o_1
X_13918_ net1071 game.CPU.applesa.ab.check_walls.above.walls\[152\] vssd1 vssd1 vccd1
+ vccd1 _07792_ sky130_fd_sc_hd__xor2_1
X_14898_ net1105 _08414_ vssd1 vssd1 vccd1 vccd1 _08675_ sky130_fd_sc_hd__and2_1
X_17686_ game.CPU.walls.rand_wall.count_luck\[4\] _03068_ vssd1 vssd1 vccd1 vccd1
+ _03070_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_348_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_334_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19425_ clknet_leaf_39_clk game.writer.tracker.next_frame\[20\] net1332 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[20\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19071__CLK net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13849_ game.writer.tracker.frame\[566\] net845 net708 game.writer.tracker.frame\[567\]
+ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__o22a_1
X_16637_ net118 _02536_ net557 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_256_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_231_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18639__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19356_ clknet_leaf_71_clk game.CPU.applesa.twoapples.absxs.next_head\[1\] vssd1
+ vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.x_final\[1\] sky130_fd_sc_hd__dfxtp_1
X_16568_ net1634 _02488_ _02492_ net127 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[86\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19189__D net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11598__A2 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18307_ net641 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
X_15519_ net853 net841 net859 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16499_ _02290_ net235 net206 net198 vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__and4b_4
X_19287_ clknet_leaf_69_clk net405 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.y_final\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_98_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13419__S0 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09040_ game.CPU.applesa.ab.absxs.body_x\[11\] vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__inv_2
XFILLER_0_304_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15733__A1 game.CPU.applesa.ab.absxs.body_y\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18238_ net665 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XFILLER_0_303_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16930__B1 _02650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12208__B net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18789__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11112__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_288_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09412__A1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18169_ net629 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__inv_2
XANTENNA__09412__B2 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10558__B1 _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 _08652_ vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 game.writer.tracker.frame\[276\] vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_345_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold424 game.CPU.randy.f1.a1.count\[2\] vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 game.writer.tracker.frame\[51\] vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_269_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold446 game.writer.tracker.frame\[542\] vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload31_A clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold457 game.writer.tracker.frame\[532\] vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 game.writer.tracker.frame\[267\] vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__A3 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_267_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09942_ net1114 _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__nand2_1
Xhold479 game.writer.tracker.frame\[530\] vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 net905 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__buf_6
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_209_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout915 net918 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__buf_4
XFILLER_0_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout926 net928 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_216_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09873_ net927 game.CPU.applesa.ab.absxs.body_x\[111\] game.CPU.applesa.ab.absxs.body_x\[109\]
+ net917 _04110_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__a221o_1
Xfanout937 _03190_ vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__clkbuf_2
Xfanout948 net950 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout294_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19731__RESET_B net1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 net982 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1001_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16461__A2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_224_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09533__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18619__Q game.CPU.applesa.ab.absxs.body_y\[113\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19414__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout559_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_224_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_356_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12483__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13680__C1 net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout726_A _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16764__A3 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_X net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19564__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13432__C1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09307_ net904 game.CPU.applesa.ab.absxs.body_y\[54\] _03308_ net1159 vssd1 vssd1
+ vccd1 vccd1 _03550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_354_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1256_X net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11303__A game.CPU.applesa.ab.apple_possible\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_106_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09238_ net780 vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__inv_2
XANTENNA__14527__A2 _08400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_302_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12538__A1 game.CPU.applesa.ab.absxs.body_x\[40\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11022__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ game.CPU.applesa.ab.check_walls.above.walls\[68\] vssd1 vssd1 vccd1 vccd1
+ _03418_ sky130_fd_sc_hd__inv_2
XANTENNA__09403__A1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09403__B2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11200_ game.CPU.applesa.ab.absxs.body_x\[23\] net544 net538 game.CPU.applesa.ab.absxs.body_y\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09708__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_309_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12180_ _06004_ _06034_ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14333__B net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19819__RESET_B net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ _03303_ net401 vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09427__B game.CPU.applesa.ab.check_walls.above.walls\[113\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15148__C game.CPU.applesa.ab.check_walls.above.walls\[176\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12134__A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17229__A1 _02412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14160__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11062_ game.CPU.applesa.ab.absxs.body_y\[24\] net533 vssd1 vssd1 vccd1 vccd1 _04952_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_247_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13664__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13517__X _07391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ net1153 _04220_ _04219_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__a21boi_1
XANTENNA__11973__A game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15870_ _03281_ net269 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10721__B1 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19401__RESET_B net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16452__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ _08626_ _08627_ vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__nor2_1
XANTENNA__09443__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_240_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17540_ _04808_ _02818_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__and2b_1
X_14752_ game.CPU.randy.counter1.count1\[16\] _08573_ vssd1 vssd1 vccd1 vccd1 _08576_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_263_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11964_ _05844_ _05851_ _05819_ _05830_ _05843_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_203_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19907__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13703_ game.writer.tracker.frame\[501\] game.writer.tracker.frame\[503\] game.writer.tracker.frame\[504\]
+ game.writer.tracker.frame\[502\] net975 net1015 vssd1 vssd1 vccd1 vccd1 _07577_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10915_ net414 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.next_head\[1\] sky130_fd_sc_hd__inv_2
XFILLER_0_86_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17471_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14683_ _08518_ _08520_ _08521_ _08505_ vssd1 vssd1 vccd1 vccd1 _08522_ sky130_fd_sc_hd__a31o_1
XANTENNA__16276__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_230_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11895_ net821 net303 vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__nand2_1
XFILLER_0_183_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19210_ net1167 _00022_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_possible\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13634_ _07506_ _07507_ net495 vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__mux2_1
X_16422_ net134 net114 _02372_ _02387_ net725 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__o41a_2
XFILLER_0_128_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10846_ _03506_ game.CPU.randy.counter1.count1\[7\] _03507_ game.CPU.randy.counter1.count1\[6\]
+ _04748_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14508__B net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16353_ game.writer.tracker.frame\[26\] net734 _02337_ vssd1 vssd1 vccd1 vccd1 _02338_
+ sky130_fd_sc_hd__and3_1
X_19141_ net1184 _00183_ _00812_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[186\]
+ sky130_fd_sc_hd__dfrtp_4
X_13565_ game.writer.tracker.frame\[361\] game.writer.tracker.frame\[363\] game.writer.tracker.frame\[364\]
+ game.writer.tracker.frame\[362\] net968 net1001 vssd1 vssd1 vccd1 vccd1 _07439_
+ sky130_fd_sc_hd__mux4_1
X_10777_ net933 game.CPU.applesa.ab.absxs.body_y\[55\] vssd1 vssd1 vccd1 vccd1 _04720_
+ sky130_fd_sc_hd__and2_1
XANTENNA__18931__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15304_ game.CPU.applesa.twomode.number\[6\] _08846_ game.CPU.applesa.twomode.counter
+ vssd1 vssd1 vccd1 vccd1 _08852_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12516_ game.CPU.applesa.ab.absxs.body_y\[68\] net362 vssd1 vssd1 vccd1 vccd1 _06393_
+ sky130_fd_sc_hd__xnor2_1
X_19072_ net1185 _00107_ _00743_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_325_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16284_ net70 _02286_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13496_ _07063_ _07078_ net689 vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17180__A3 _02479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13726__B1 _07599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13839__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18023_ net662 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__inv_2
X_15235_ game.CPU.applesa.normal1.number\[3\] _08795_ vssd1 vssd1 vccd1 vccd1 _08798_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_251_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12447_ game.CPU.applesa.ab.absxs.body_y\[91\] net364 vssd1 vssd1 vccd1 vccd1 _06324_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_301_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14524__A _07164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap357_A _08416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_288_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15166_ net1226 net1253 game.CPU.walls.rand_wall.x_final\[2\] vssd1 vssd1 vccd1 vccd1
+ _00210_ sky130_fd_sc_hd__and3_1
XANTENNA__09618__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12378_ _03322_ game.CPU.applesa.twoapples.absxs.next_head\[6\] net366 game.CPU.applesa.ab.absxs.body_y\[115\]
+ _06254_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__o221a_1
XANTENNA__19095__Q game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14117_ game.CPU.applesa.ab.check_walls.above.walls\[173\] net862 net1052 _03471_
+ vssd1 vssd1 vccd1 vccd1 _07991_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_22_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11329_ game.CPU.applesa.ab.check_walls.above.walls\[85\] net314 vssd1 vssd1 vccd1
+ vccd1 _05218_ sky130_fd_sc_hd__and2_1
X_19974_ clknet_leaf_39_clk game.writer.tracker.next_frame\[569\] net1331 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[569\] sky130_fd_sc_hd__dfrtp_1
X_15097_ net1203 net1229 net795 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14151__B1 _07766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16691__A2 _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14048_ net1043 game.CPU.applesa.ab.check_walls.above.walls\[195\] vssd1 vssd1 vccd1
+ vccd1 _07922_ sky130_fd_sc_hd__xor2_1
X_18925_ clknet_leaf_5_clk net1393 _00609_ vssd1 vssd1 vccd1 vccd1 game.CPU.left_button.eD1.D
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_253_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19437__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13574__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11883__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_340_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18856_ clknet_leaf_0_clk _01247_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16979__B1 _02665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17807_ net944 _03139_ _03140_ _03142_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__a22o_1
XFILLER_0_206_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15074__B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18787_ clknet_leaf_3_clk game.CPU.state1.Qn\[1\] _00524_ vssd1 vssd1 vccd1 vccd1
+ game.CPU.clock1.game_state\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10499__A _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15999_ game.CPU.applesa.ab.check_walls.above.walls\[97\] net472 net458 game.CPU.applesa.ab.check_walls.above.walls\[99\]
+ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__o22a_1
X_17738_ game.CPU.applesa.ab.count\[2\] game.CPU.applesa.ab.count\[1\] game.CPU.applesa.ab.count\[3\]
+ _03101_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__nand4_2
XANTENNA__19587__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11107__B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17669_ game.CPU.kyle.L1.cnt_500hz\[12\] game.CPU.kyle.L1.cnt_500hz\[13\] _03053_
+ game.CPU.kyle.L1.cnt_500hz\[14\] vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_11_Left_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15090__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19408_ clknet_leaf_48_clk game.writer.tracker.next_frame\[3\] net1295 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14418__B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10946__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13965__B1 game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19339_ clknet_leaf_72_clk _01355_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.count_luck\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09633__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_351_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12219__A _03381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09633__B2 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11123__A game.CPU.applesa.ab.absxs.body_y\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10243__A2 game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_289_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13749__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09023_ game.CPU.applesa.ab.absxs.body_x\[50\] vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13812__S0 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout307_A _05606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1049_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold210 game.writer.tracker.frame\[506\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19983__RESET_B net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09528__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14390__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold221 game.writer.tracker.frame\[348\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11777__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold232 game.writer.tracker.frame\[309\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_276_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_269_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold243 game.writer.tracker.frame\[548\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 game.writer.tracker.frame\[323\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19912__RESET_B net1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold265 game.writer.tracker.frame\[465\] vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold276 game.writer.tracker.frame\[210\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 game.writer.tracker.frame\[186\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1216_A game.CPU.walls.rand_wall.start_enable vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10951__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout701 net707 vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_284_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout712 _06594_ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_2
Xhold298 game.writer.tracker.frame\[42\] vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14142__B1 _07983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09925_ net1092 net847 _04165_ vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__a21o_1
Xfanout723 net724 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_187_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout734 net738 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_2
XANTENNA_fanout676_A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 _04451_ vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__clkbuf_4
X_20045_ game.dcx vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_2
X_09856_ net1131 game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1 _04099_
+ sky130_fd_sc_hd__or2_1
Xfanout767 game.CPU.applesa.ab.apple_possible\[2\] vssd1 vssd1 vccd1 vccd1 net767
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_129_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_304_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1004_X net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout778 net779 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__buf_4
XANTENNA__10703__B1 _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18804__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout789 game.CPU.applesa.ab.check_walls.above.walls\[151\] vssd1 vssd1 vccd1 vccd1
+ net789 sky130_fd_sc_hd__buf_2
XFILLER_0_213_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09787_ _04022_ _04023_ _04028_ _04029_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout843_A _06574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12401__B net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16985__A3 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12456__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10202__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_202_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15712__B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_276_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09872__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18954__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09872__B2 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ game.CPU.applesa.ab.absxs.body_y\[78\] _04623_ _04624_ game.CPU.applesa.ab.absxs.body_y\[74\]
+ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ game.CPU.applesa.ab.check_walls.above.walls\[59\] net764 vssd1 vssd1 vccd1
+ vccd1 _05569_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_138_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_327_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14328__B net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ _04683_ game.CPU.applesa.ab.absxs.body_x\[57\] net327 vssd1 vssd1 vccd1 vccd1
+ _01120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_342_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_313_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12129__A game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16824__A net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13800__X _07674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12854__S1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_180_Left_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13350_ net213 _07222_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__and2_1
XFILLER_0_307_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10562_ net1123 _04156_ _04645_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_8_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17162__A3 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13708__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12301_ game.CPU.applesa.ab.check_walls.above.walls\[45\] net549 vssd1 vssd1 vccd1
+ vccd1 _06187_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11968__A game.CPU.applesa.ab.check_walls.above.walls\[148\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ game.writer.tracker.frame\[458\] game.writer.tracker.frame\[459\] net1011
+ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__mux2_1
X_10493_ _04608_ _04613_ _04614_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09388__B1 game.CPU.applesa.ab.check_walls.above.walls\[165\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15020_ net1228 net1256 game.CPU.applesa.ab.check_walls.above.walls\[48\] vssd1 vssd1
+ vccd1 vccd1 _00239_ sky130_fd_sc_hd__and3_1
XFILLER_0_267_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14381__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12232_ _06117_ _06023_ _06022_ _06116_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_279_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15159__B net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_287_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19653__RESET_B net1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ _05524_ _05528_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__nand2_1
XFILLER_0_248_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_229_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14998__B net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11114_ _04994_ _04995_ _04997_ _04998_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a22o_1
X_16971_ _02436_ net96 _02661_ game.writer.tracker.frame\[320\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[320\] sky130_fd_sc_hd__a22o_1
XFILLER_0_275_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12094_ _05489_ _05490_ _05492_ _05495_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__or4b_1
XANTENNA__13394__S net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18710_ clknet_leaf_52_clk _01127_ _00447_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[72\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11498__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11045_ game.CPU.applesa.ab.absxs.body_x\[83\] net546 vssd1 vssd1 vccd1 vccd1 _04935_
+ sky130_fd_sc_hd__xnor2_1
X_15922_ game.CPU.applesa.ab.check_walls.above.walls\[135\] net430 vssd1 vssd1 vccd1
+ vccd1 _01934_ sky130_fd_sc_hd__xnor2_1
X_19690_ clknet_leaf_34_clk game.writer.tracker.next_frame\[285\] net1313 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[285\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16425__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18641_ clknet_leaf_59_clk _01058_ _00378_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[39\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_265_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10077__C_N _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15853_ game.CPU.applesa.ab.absxs.body_y\[98\] _08429_ vssd1 vssd1 vccd1 vccd1 _01865_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_204_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12311__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14804_ game.CPU.randy.counter1.count\[9\] _08614_ net138 vssd1 vssd1 vccd1 vccd1
+ _08617_ sky130_fd_sc_hd__o21ai_1
X_18572_ clknet_leaf_62_clk _00992_ _00309_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_12996_ game.writer.tracker.frame\[522\] game.writer.tracker.frame\[523\] net1004
+ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__mux2_1
X_15784_ _03332_ net339 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16718__B _02289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17523_ _02950_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__inv_2
XANTENNA__15622__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11947_ game.CPU.applesa.ab.check_walls.above.walls\[118\] net299 vssd1 vssd1 vccd1
+ vccd1 _05835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14735_ net55 _08563_ _08564_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__and3_1
XANTENNA__16189__B2 game.CPU.applesa.ab.absxs.body_y\[69\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09863__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14519__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__B2 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16728__A3 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_345_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_290_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11670__A1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17454_ net1121 _02786_ _02882_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__o21a_1
X_14666_ game.CPU.randy.counter1.count1\[8\] _08504_ vssd1 vssd1 vccd1 vccd1 _08505_
+ sky130_fd_sc_hd__and2_1
X_11878_ net569 _05236_ _05241_ _05242_ _05765_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__o2111a_1
XANTENNA__11670__B2 game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_253_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14238__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13617_ _07489_ _07490_ net515 vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__mux2_1
X_16405_ net1793 _02371_ _02375_ net111 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[40\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10829_ _04482_ _04567_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__or2_2
XFILLER_0_144_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17138__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14597_ game.CPU.clock1.counter\[3\] _08455_ net739 vssd1 vssd1 vccd1 vccd1 _08456_
+ sky130_fd_sc_hd__a21oi_1
X_17385_ net1124 _02785_ _02811_ _02814_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__a211o_1
XFILLER_0_223_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19124_ net1183 _00164_ _00795_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[169\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_144_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16336_ net225 _02326_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__nor2_8
X_13548_ game.writer.tracker.frame\[73\] game.writer.tracker.frame\[75\] game.writer.tracker.frame\[76\]
+ game.writer.tracker.frame\[74\] net974 net1010 vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_298_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18722__Q game.CPU.applesa.ab.absxs.body_x\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16267_ _02236_ _02271_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__nor2_8
X_19055_ net1192 _00089_ _00726_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[100\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13479_ net487 _07350_ _07352_ net209 vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_329_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16900__A3 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15218_ game.CPU.applesa.normal1.number\[4\] _08778_ vssd1 vssd1 vccd1 vccd1 _08784_
+ sky130_fd_sc_hd__nand2_1
X_18006_ net613 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
XFILLER_0_298_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_258_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14372__B1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09348__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16198_ _01627_ _01632_ _02208_ _02209_ _02121_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__o32a_1
XANTENNA__19394__RESET_B net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15149_ net1213 net1239 game.CPU.applesa.ab.check_walls.above.walls\[177\] vssd1
+ vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_266_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18827__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_264_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_318_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19957_ clknet_leaf_43_clk game.writer.tracker.next_frame\[552\] net1305 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[552\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_206_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10006__B _04212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ net922 game.CPU.applesa.ab.absxs.body_x\[22\] game.CPU.applesa.ab.absxs.body_y\[21\]
+ net900 _03951_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__a221o_1
XANTENNA__15085__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18908_ clknet_leaf_4_clk _01275_ _00592_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[6\]
+ sky130_fd_sc_hd__dfstp_4
X_19888_ clknet_leaf_27_clk game.writer.tracker.next_frame\[483\] net1309 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[483\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_254_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16416__A2 _02299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ net1127 net788 vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_6_clk_X clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18839_ clknet_leaf_73_clk _01230_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_334_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12438__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ _03808_ _03809_ _03810_ _03814_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_353_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09811__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14429__A game.CPU.applesa.ab.absxs.body_y\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout257_A _05207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11661__A1 game.CPU.applesa.ab.check_walls.above.walls\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10464__A2 game.CPU.applesa.ab.absxs.body_x\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10676__B _04701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_186_Right_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16644__A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17459__B _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16363__B net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17144__A3 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11788__A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18632__Q game.CPU.applesa.ab.absxs.body_y\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19602__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12236__X _06122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1333_A net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09006_ game.CPU.applesa.ab.absxs.body_x\[104\] vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_189_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14363__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_276_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_306_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19752__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15707__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout960_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 net522 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_4
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout531 net532 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__buf_4
Xfanout542 net543 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_8
X_09908_ net1109 _04148_ _04149_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__nand3_1
XFILLER_0_272_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__clkbuf_4
Xfanout564 net565 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_4
XFILLER_0_272_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout575 _04443_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09542__B1 game.CPU.applesa.ab.XMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout586 net587 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__buf_4
X_09839_ net904 game.CPU.applesa.ab.absxs.body_y\[106\] _03321_ net1159 vssd1 vssd1
+ vccd1 vccd1 _04082_ sky130_fd_sc_hd__o22a_1
Xfanout597 net598 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_4
X_20028_ net1276 vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_272_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout846_X net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_244_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16958__A3 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ game.writer.tracker.frame\[272\] game.writer.tracker.frame\[273\] net1001
+ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__mux2_2
XFILLER_0_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15723__A game.CPU.applesa.ab.absxs.body_y\[52\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16538__B net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11801_ _05680_ _05681_ _05688_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__or3_2
XFILLER_0_96_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_347_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_317_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ game.writer.tracker.frame\[92\] game.writer.tracker.frame\[93\] net1019 vssd1
+ vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__mux2_1
X_14520_ _08393_ vssd1 vssd1 vccd1 vccd1 _08394_ sky130_fd_sc_hd__inv_2
XANTENNA__19132__CLK net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11732_ net749 _05478_ _05476_ net570 vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11652__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11652__B2 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14058__B game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14451_ game.CPU.applesa.ab.absxs.body_y\[14\] net953 vssd1 vssd1 vccd1 vccd1 _08325_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_354_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11663_ game.CPU.applesa.ab.check_walls.above.walls\[122\] net765 vssd1 vssd1 vccd1
+ vccd1 _05552_ sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16591__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13402_ _06865_ _06877_ net685 vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__mux2_1
X_17170_ net149 _02466_ net73 _02723_ net1523 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[457\]
+ sky130_fd_sc_hd__a32o_1
X_10614_ game.CPU.applesa.ab.absxs.body_x\[75\] _04675_ _04676_ game.CPU.applesa.ab.absxs.body_x\[71\]
+ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14382_ game.CPU.applesa.ab.absxs.body_x\[81\] net1060 vssd1 vssd1 vccd1 vccd1 _08256_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__11404__B2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_289_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11594_ net743 _05478_ _05479_ _05481_ _05477_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17135__A3 _02690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13389__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19287__D net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16121_ game.CPU.applesa.ab.check_walls.above.walls\[178\] net466 net333 _03479_
+ _02132_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a221o_2
X_13333_ net677 _06738_ _07206_ net200 vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__o211a_1
XANTENNA__19282__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10545_ _04584_ _04607_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__nor2_2
XFILLER_0_323_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09168__A game.CPU.applesa.ab.check_walls.above.walls\[67\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14354__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16052_ _03294_ net339 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__xnor2_1
X_13264_ net502 _07135_ _07137_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__a21o_1
X_10476_ game.CPU.applesa.ab.absxs.body_x\[93\] _04601_ _04604_ net929 vssd1 vssd1
+ vccd1 vccd1 _01196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_295_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15003_ net1223 net1251 net825 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__and3_1
X_12215_ _06097_ _06098_ _06099_ _06100_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__or4_2
XANTENNA__11210__B net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_295_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13195_ game.writer.tracker.frame\[406\] game.writer.tracker.frame\[407\] net1037
+ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19811_ clknet_leaf_39_clk game.writer.tracker.next_frame\[406\] net1353 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[406\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09781__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ net781 net295 net292 game.CPU.applesa.ab.check_walls.above.walls\[190\] vssd1
+ vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__15617__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10391__A1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10391__B2 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_285_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19742_ clknet_leaf_25_clk game.writer.tracker.next_frame\[337\] net1322 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[337\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12668__A0 game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16954_ _02408_ net94 _02657_ net1664 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[307\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09615__B game.CPU.applesa.ab.check_walls.above.walls\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12077_ net808 net293 vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__or2_1
XANTENNA__13865__C1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15905_ game.CPU.applesa.ab.absxs.body_x\[56\] net355 vssd1 vssd1 vccd1 vccd1 _01917_
+ sky130_fd_sc_hd__xnor2_1
X_11028_ game.CPU.applesa.ab.absxs.body_x\[64\] net325 vssd1 vssd1 vccd1 vccd1 _04918_
+ sky130_fd_sc_hd__nand2_1
X_19673_ clknet_leaf_30_clk game.writer.tracker.next_frame\[268\] net1285 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[268\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_288_Right_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16885_ net1797 _02631_ net93 _02452_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[259\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11583__D _05471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14409__A1 game.CPU.applesa.ab.absxs.body_x\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13880__A2 game.CPU.applesa.ab.check_walls.above.walls\[106\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17071__A2 net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18624_ clknet_leaf_11_clk _01041_ _00361_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[106\]
+ sky130_fd_sc_hd__dfrtp_4
X_15836_ _03259_ net351 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11891__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11055__A1_N game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09631__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18555_ clknet_leaf_45_clk _00978_ net1279 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.cmd_num\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12979_ net219 _06606_ net282 vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__a21o_1
XANTENNA__09836__A1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15767_ game.CPU.applesa.ab.absxs.body_x\[116\] net355 net452 game.CPU.applesa.ab.absxs.body_y\[116\]
+ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13632__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_304_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09836__B2 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17506_ _02927_ _02931_ _02932_ _02934_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__or4_1
XFILLER_0_318_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14718_ game.CPU.randy.counter1.count1\[5\] game.CPU.randy.counter1.count1\[4\] _08548_
+ vssd1 vssd1 vccd1 vccd1 _08553_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18486_ net630 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15698_ game.CPU.applesa.ab.absxs.body_x\[31\] net457 net438 game.CPU.applesa.ab.absxs.body_y\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_43_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17437_ _02844_ _02858_ _02860_ _02866_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__or4_1
XANTENNA__19625__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14649_ game.CPU.randy.f1.state\[3\] game.CPU.randy.f1.state\[2\] game.CPU.randy.f1.state\[0\]
+ game.CPU.randy.f1.state\[1\] vssd1 vssd1 vccd1 vccd1 _08488_ sky130_fd_sc_hd__or4b_1
XANTENNA_16 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_311_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_27 _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13396__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_38 game.writer.tracker.frame\[336\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_49 game.writer.tracker.frame\[305\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17368_ _08748_ _02788_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__or2_1
XANTENNA__17126__A3 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19575__RESET_B net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19107_ net1180 _00146_ _00778_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[152\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_314_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16319_ _02245_ net235 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17299_ net1975 net722 _02756_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[553\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__13148__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19775__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19038_ net1193 _00269_ _00709_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[83\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14345__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_212_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12216__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11120__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10017__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16098__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09365__X _03608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__A1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19005__CLK net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__B2 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12659__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13856__C1 net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13320__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12123__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_254_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_301_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_255_Right_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16198__X _02210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_345_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13871__A2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ net1103 game.CPU.applesa.ab.check_walls.above.walls\[1\] vssd1 vssd1 vccd1
+ vccd1 _03867_ sky130_fd_sc_hd__xor2_1
XFILLER_0_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17062__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19155__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16358__B _02301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09555_ net1094 game.CPU.applesa.ab.absxs.body_x\[62\] vssd1 vssd1 vccd1 vccd1 _03798_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__13084__B1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout162_X net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1283_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout639_A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10437__A2 _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ net920 game.CPU.applesa.ab.check_walls.above.walls\[186\] _03483_ net1135
+ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_273_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_336_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_352_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1071_X net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16573__B2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_A game.CPU.applesa.ab.check_walls.above.walls\[93\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_X net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_351_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_312_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16093__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_305_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11311__A game.CPU.applesa.ab.check_walls.above.walls\[65\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10330_ net740 _04488_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__nand2_1
XANTENNA__16876__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13234__S1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_249_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_239_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11030__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12898__A0 _06768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ _04452_ _04453_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_284_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12000_ game.CPU.applesa.ab.check_walls.above.walls\[165\] net386 vssd1 vssd1 vccd1
+ vccd1 _05887_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_226_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10192_ net1097 _04383_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout963_X net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1304 net1305 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__clkbuf_4
Xfanout1315 net1316 vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_319_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1326 net1327 vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__clkbuf_4
Xfanout1337 net1359 vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__clkbuf_4
Xfanout1348 net1359 vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__clkbuf_4
Xfanout350 net353 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_148_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout75_X net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout361 net362 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_323_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1359 net1360 vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13311__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout372 net374 vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_4
XFILLER_0_260_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout383 net384 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_2
XANTENNA__10125__A1 net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13951_ net867 net793 _03450_ net947 vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout394 net395 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13862__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13525__X _07399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_222_Right_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12902_ game.writer.tracker.frame\[18\] game.writer.tracker.frame\[19\] net1024 vssd1
+ vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__mux2_1
X_16670_ net168 net154 net56 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__and3_1
X_13882_ net963 game.CPU.applesa.ab.check_walls.above.walls\[101\] vssd1 vssd1 vccd1
+ vccd1 _07756_ sky130_fd_sc_hd__xor2_1
XANTENNA__16800__A2 _02322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12833_ game.writer.tracker.frame\[286\] game.writer.tracker.frame\[287\] net1012
+ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__mux2_1
X_15621_ _03423_ net270 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19648__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09818__A1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09818__B2 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_295_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16086__A1_N game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18340_ net595 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__inv_2
XFILLER_0_271_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12764_ _06632_ _06633_ _06635_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__nor4_1
X_15552_ net965 net954 net943 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_237_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16555__Y _02484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14503_ game.CPU.apple_location\[0\] net886 net852 game.CPU.apple_location\[6\] vssd1
+ vssd1 vccd1 vccd1 _08377_ sky130_fd_sc_hd__a22o_1
X_11715_ net765 net759 _04441_ game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1
+ vccd1 vccd1 _05603_ sky130_fd_sc_hd__a31o_1
X_15483_ _08927_ _08931_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__or2_2
X_18271_ net662 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11205__B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15900__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12695_ _06565_ _06567_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__xor2_2
XANTENNA__14356__X _08230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16284__A net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13378__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16715__C net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17222_ _02396_ net142 net119 _02736_ net1612 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[496\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19798__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14434_ _03351_ net984 net939 _03348_ _08302_ vssd1 vssd1 vccd1 vccd1 _08308_ sky130_fd_sc_hd__a221o_1
XANTENNA__18672__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11646_ game.CPU.applesa.ab.check_walls.above.walls\[9\] net772 vssd1 vssd1 vccd1
+ vccd1 _05535_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17108__A3 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_342_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17153_ _02431_ net58 _02717_ net1677 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[446\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09169__Y _03418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14365_ _08232_ _08236_ _08237_ _08238_ vssd1 vssd1 vccd1 vccd1 _08239_ sky130_fd_sc_hd__or4_1
X_11577_ net793 net249 _05464_ _05465_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__o211a_1
X_13316_ net510 _06719_ net703 vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__a21o_1
X_16104_ game.CPU.applesa.ab.absxs.body_x\[18\] net469 vssd1 vssd1 vccd1 vccd1 _02116_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__16867__A2 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17084_ net206 _02389_ net57 _02697_ net1815 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[397\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_268_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10528_ game.CPU.applesa.ab.absxs.body_x\[54\] _04609_ _04637_ game.CPU.applesa.ab.absxs.body_x\[50\]
+ vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_311_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14296_ game.CPU.applesa.ab.absxs.body_x\[53\] net1067 vssd1 vssd1 vccd1 vccd1 _08170_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_357_Right_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_326_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13247_ net209 _07120_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__or2_1
XFILLER_0_295_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16035_ game.CPU.applesa.ab.absxs.body_y\[47\] net434 vssd1 vssd1 vccd1 vccd1 _02047_
+ sky130_fd_sc_hd__nor2_1
X_10459_ _04589_ _04593_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__and2_4
XANTENNA__18004__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_248_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16619__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09626__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ _07048_ _07049_ _07050_ _07051_ net499 net689 vssd1 vssd1 vccd1 vccd1 _07052_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_283_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11875__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_261_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12129_ game.CPU.applesa.ab.check_walls.above.walls\[5\] net389 vssd1 vssd1 vccd1
+ vccd1 _06016_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_229_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19178__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__B game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17986_ net614 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__inv_2
XANTENNA__15066__C game.CPU.applesa.ab.check_walls.above.walls\[94\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13302__A1 _06768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19725_ clknet_leaf_35_clk game.writer.tracker.next_frame\[320\] net1346 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[320\] sky130_fd_sc_hd__dfrtp_1
X_16937_ net163 net68 net87 _02652_ net1560 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[295\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__10116__A1 game.CPU.applesa.enable_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16459__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_251_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17044__A2 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19656_ clknet_leaf_23_clk game.writer.tracker.next_frame\[251\] net1348 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[251\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10667__A2 _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16868_ net153 _02423_ net107 _02628_ net1541 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[250\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_315_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_337_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18607_ clknet_leaf_69_clk _01024_ _00344_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[89\]
+ sky130_fd_sc_hd__dfrtp_4
X_15819_ game.CPU.applesa.ab.absxs.body_x\[90\] net465 vssd1 vssd1 vccd1 vccd1 _01831_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__15082__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19587_ clknet_leaf_36_clk game.writer.tracker.next_frame\[182\] net1351 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[182\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09809__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16799_ _02483_ net103 _02600_ game.writer.tracker.frame\[209\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[209\] sky130_fd_sc_hd__a22o_1
XFILLER_0_87_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09809__B2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09340_ game.CPU.applesa.ab.absxs.body_y\[89\] net898 net1107 _03264_ vssd1 vssd1
+ vccd1 vccd1 _03583_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_259_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18538_ net611 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16465__Y _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09271_ game.CPU.clock1.counter\[6\] vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__inv_2
XFILLER_0_334_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18469_ net652 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__inv_2
XANTENNA__15810__B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_306_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload61_A clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11919__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout122_A _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14318__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16858__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_348_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_324_Right_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1031_A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17807__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09745__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11785__B net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17283__A2 _02577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_299_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08986_ game.CPU.applesa.ab.absxs.body_x\[79\] vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__inv_2
XFILLER_0_199_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_270_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19741__Q game.writer.tracker.frame\[336\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16369__A _06573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17035__A2 _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10658__A2 _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Left_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_197_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09607_ net1085 _03285_ _03355_ net1159 vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout923_A _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__A game.CPU.applesa.ab.apple_possible\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12804__A0 game.writer.tracker.frame\[336\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11607__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ net1137 net812 vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__xor2_1
XANTENNA__18695__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16375__Y _02354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19940__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11025__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_241_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15720__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09469_ net1083 _03228_ game.CPU.applesa.ab.absxs.body_x\[94\] net921 _03708_ vssd1
+ vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__a221o_1
X_11500_ net746 _05385_ _05388_ net564 vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__o22a_1
XFILLER_0_171_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14557__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12480_ game.CPU.applesa.ab.absxs.body_y\[30\] net517 net370 game.CPU.applesa.ab.absxs.body_x\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19188__Q game.CPU.walls.rand_wall.start_enable vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ game.CPU.applesa.ab.check_walls.above.walls\[24\] net777 vssd1 vssd1 vccd1
+ vccd1 _05320_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_321_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_232_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14150_ _07882_ _07884_ _07755_ vssd1 vssd1 vccd1 vccd1 _08024_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_34_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16849__A2 _02391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11362_ net824 net252 net317 net823 vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__o22a_1
X_13101_ net491 _06974_ _06973_ net228 vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__o211a_1
XANTENNA__10594__B2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11976__A game.CPU.applesa.ab.apple_possible\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10313_ game.CPU.randy.f1.a1.count\[14\] _04495_ vssd1 vssd1 vccd1 vccd1 _04496_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__15448__A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14081_ net1046 game.CPU.applesa.ab.check_walls.above.walls\[91\] vssd1 vssd1 vccd1
+ vccd1 _07955_ sky130_fd_sc_hd__xor2_1
XANTENNA__10880__A game.CPU.applesa.ab.apple_possible\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11293_ _04908_ _04909_ _04915_ _04916_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__a22o_1
XANTENNA__14352__A game.CPU.applesa.ab.absxs.body_x\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13032_ net680 _06890_ _06905_ net507 vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__o211a_1
XANTENNA__19320__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09736__B1 game.CPU.applesa.ab.absxs.body_y\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11695__B net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ game.CPU.applesa.ab.count_luck\[4\] game.CPU.applesa.ab.count_luck\[5\] game.CPU.applesa.ab.count_luck\[1\]
+ _04422_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__a31o_1
XFILLER_0_266_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14071__B game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1101 game.CPU.applesa.ab.snake_head_x\[1\] vssd1 vssd1 vccd1 vccd1 net1101
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA__17274__A2 _02258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17840_ _03166_ _03167_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__nor2_1
Xfanout1112 net1113 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10175_ net897 _04367_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1123 game.CPU.bodymain1.main.score\[1\] vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_31_clk_X clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1134 net1135 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__buf_4
Xfanout1145 net1152 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__buf_4
Xfanout1156 net1157 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__clkbuf_2
Xfanout1167 net1169 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__buf_2
X_17771_ game.CPU.applesa.twoapples.count_luck\[6\] _03121_ game.CPU.applesa.twoapples.count_luck\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__a21o_1
XFILLER_0_273_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14983_ net1227 net1252 game.CPU.applesa.ab.check_walls.above.walls\[11\] vssd1 vssd1
+ vccd1 vccd1 _00198_ sky130_fd_sc_hd__and3_1
XANTENNA__19470__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16279__A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_233_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1178 net1179 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_233_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19510_ clknet_leaf_14_clk game.writer.tracker.next_frame\[105\] net1282 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[105\] sky130_fd_sc_hd__dfrtp_1
Xfanout191 _06588_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_4
Xfanout1189 net1190 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__buf_2
X_16722_ net1970 _02575_ _02576_ net106 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[156\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13391__S0 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17026__A2 _02670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11846__A1 game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13934_ net890 game.CPU.applesa.ab.check_walls.above.walls\[32\] net824 net869 vssd1
+ vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09181__A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19441_ clknet_leaf_43_clk game.writer.tracker.next_frame\[36\] net1299 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[36\] sky130_fd_sc_hd__dfrtp_1
X_16653_ net1952 _02543_ _02544_ net128 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[119\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13048__B1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16785__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13865_ net240 _07735_ _07738_ _07730_ net207 vssd1 vssd1 vccd1 vccd1 _07739_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_18_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16566__X _02491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_46_clk_X clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18494__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_347_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15604_ game.CPU.applesa.ab.check_walls.above.walls\[115\] net457 net332 _03442_
+ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__a22o_1
X_12816_ game.writer.tracker.frame\[328\] game.writer.tracker.frame\[329\] net1015
+ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__mux2_2
XFILLER_0_186_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19372_ clknet_leaf_70_clk _01378_ _00953_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location2\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12105__A2_N net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16584_ _02427_ net144 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_158_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13796_ game.writer.tracker.frame\[390\] net843 net674 game.writer.tracker.frame\[392\]
+ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__o22a_1
XFILLER_0_84_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14260__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18323_ net615 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
X_15535_ _01523_ _01546_ _01507_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_316_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12747_ game.writer.tracker.frame\[76\] game.writer.tracker.frame\[77\] net999 vssd1
+ vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__mux2_1
XANTENNA__16537__B2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13431__A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_315_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18254_ net644 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
X_15466_ game.writer.updater.commands.count\[7\] game.writer.updater.commands.count\[6\]
+ game.writer.updater.commands.count\[5\] vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__and3_1
X_12678_ net1057 net1048 vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_332_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19098__Q game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14246__B net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17205_ _02609_ net120 _02732_ net1686 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[483\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_170_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_331_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14417_ game.CPU.applesa.ab.absxs.body_y\[109\] net964 vssd1 vssd1 vccd1 vccd1 _08291_
+ sky130_fd_sc_hd__xnor2_1
X_11629_ _05506_ _05514_ _05516_ _05517_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__or4_1
X_18185_ net609 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__inv_2
XFILLER_0_315_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15397_ _08935_ _08938_ vssd1 vssd1 vccd1 vccd1 _08939_ sky130_fd_sc_hd__or2_1
XFILLER_0_231_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17136_ _02398_ net60 _02713_ net1863 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[433\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12574__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14348_ game.CPU.applesa.ab.absxs.body_x\[34\] net1054 vssd1 vssd1 vccd1 vccd1 _08222_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10585__A1 game.CPU.applesa.ab.absxs.body_x\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold606 game.CPU.applesa.twoapples.count\[1\] vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 game.writer.tracker.frame\[572\] vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11782__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13577__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold628 game.writer.tracker.frame\[73\] vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18730__Q game.CPU.applesa.ab.absxs.body_x\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17067_ _02240_ net120 vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__nand2_1
XANTENNA__12334__X _06214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14279_ _03232_ net1053 net861 game.CPU.applesa.ab.absxs.body_y\[85\] vssd1 vssd1
+ vccd1 vccd1 _08153_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_78 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold639 game.CPU.kyle.L1.currentState\[4\] vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_268_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13523__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_256_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16018_ game.CPU.applesa.ab.absxs.body_y\[36\] net454 vssd1 vssd1 vccd1 vccd1 _02030_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_wire178_X net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15077__B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18568__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19813__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17265__A2 _02477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14079__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16473__B1 _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_326_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ net663 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__inv_2
XANTENNA__15805__B game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17017__A2 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19708_ clknet_leaf_31_clk game.writer.tracker.next_frame\[303\] net1281 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[303\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12510__A game.CPU.applesa.ab.absxs.body_x\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_224_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09342__A1_N net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19963__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19639_ clknet_leaf_28_clk game.writer.tracker.next_frame\[234\] net1290 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[234\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16776__A1 _02436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_342_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10030__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14251__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16636__B _02535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09323_ _03555_ _03561_ _03562_ _03565_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_270_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_179_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout337_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1079_A game.CPU.bad_collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ game.CPU.randy.counter1.count1\[11\] vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_192_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14156__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13437__S1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14256__A2_N net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09185_ net803 vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout504_A net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16652__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout125_X net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1246_A net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13762__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19343__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18640__Q game.CPU.applesa.ab.absxs.body_y\[38\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1034_X net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13514__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_281_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10328__B2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19493__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12404__B net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17256__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1201_X net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15715__B net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08969_ net1258 vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_145_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17008__A2 _02638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_215_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11980_ game.CPU.applesa.ab.check_walls.above.walls\[151\] net293 _05865_ _05866_
+ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__o211a_1
XANTENNA__09713__B game.CPU.applesa.ab.absxs.body_x\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_203_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10931_ game.CPU.applesa.ab.absxs.body_x\[8\] net325 vssd1 vssd1 vccd1 vccd1 _04821_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_230_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16767__A1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16386__X _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15731__A game.CPU.applesa.ab.absxs.body_x\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13650_ net279 _07513_ _07522_ _07523_ net242 vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__a221o_1
X_10862_ _04763_ _04764_ _04758_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_292_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16546__B _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12601_ _06337_ _06475_ _06476_ _06477_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__or4b_1
X_13581_ game.writer.tracker.frame\[369\] game.writer.tracker.frame\[371\] game.writer.tracker.frame\[372\]
+ game.writer.tracker.frame\[370\] net976 net1012 vssd1 vssd1 vccd1 vccd1 _07455_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__15450__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_234_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10793_ net1079 _04690_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14347__A game.CPU.applesa.ab.absxs.body_y\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_109_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15320_ game.CPU.applesa.twomode.number\[5\] _08859_ vssd1 vssd1 vccd1 vccd1 _08865_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12532_ game.CPU.applesa.ab.absxs.body_x\[98\] net370 net518 game.CPU.applesa.ab.absxs.body_y\[98\]
+ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_325_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10803__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14066__B game.CPU.applesa.ab.check_walls.above.walls\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_57_Left_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12463_ game.CPU.applesa.ab.absxs.body_y\[13\] net524 vssd1 vssd1 vccd1 vccd1 _06340_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12005__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15251_ game.CPU.kyle.L1.nextState\[5\] _08809_ net264 net1790 vssd1 vssd1 vccd1
+ vccd1 _08812_ sky130_fd_sc_hd__a22oi_4
XANTENNA__12005__B2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14202_ game.CPU.applesa.ab.absxs.body_x\[65\] net1068 vssd1 vssd1 vccd1 vccd1 _08076_
+ sky130_fd_sc_hd__xor2_1
X_11414_ net566 _05301_ _05302_ net743 vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__o22ai_1
X_15182_ _04628_ _08757_ _08755_ vssd1 vssd1 vccd1 vccd1 _08758_ sky130_fd_sc_hd__a21oi_1
X_12394_ _06262_ _06264_ _06268_ _06269_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__or4_1
XANTENNA__10567__A1 game.CPU.applesa.ab.absxs.body_x\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_73_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19646__Q game.writer.tracker.frame\[241\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10567__B2 game.CPU.applesa.ab.absxs.body_x\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14133_ net950 game.CPU.applesa.ab.check_walls.above.walls\[46\] vssd1 vssd1 vccd1
+ vccd1 _08007_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11345_ net809 net255 _05222_ _05233_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__a211o_1
XANTENNA__19836__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19990_ clknet_leaf_44_clk _01414_ net1304 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_104_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13505__A1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14064_ _07931_ _07935_ _07936_ _07937_ vssd1 vssd1 vccd1 vccd1 _07938_ sky130_fd_sc_hd__or4_1
X_18941_ net1175 _00080_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number_out\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11276_ game.CPU.applesa.ab.absxs.body_x\[62\] net409 net399 net1270 _05165_ vssd1
+ vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_37_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_245_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13015_ game.writer.tracker.frame\[540\] game.writer.tracker.frame\[541\] net1020
+ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__mux2_1
XANTENNA__17247__A2 _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ game.CPU.applesa.ab.count_luck\[1\] game.CPU.applesa.ab.count_luck\[0\] game.CPU.applesa.ab.count_luck\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__a21o_1
XANTENNA__17393__A game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18872_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[2\] _00567_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_265_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18860__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_66_Left_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19986__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17823_ game.writer.updater.commands.count\[2\] _03152_ _03154_ _03146_ vssd1 vssd1
+ vccd1 vccd1 _01411_ sky130_fd_sc_hd__o22a_1
XFILLER_0_246_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15625__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ game.CPU.randy.f1.state\[3\] game.CPU.randy.f1.state\[2\] vssd1 vssd1 vccd1
+ vccd1 _04353_ sky130_fd_sc_hd__nand2_1
XANTENNA__13269__B1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 game.CPU.start_pause_button1.sync1.Q vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_293_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17754_ game.CPU.applesa.twoapples.count_luck\[1\] _03110_ _03109_ vssd1 vssd1 vccd1
+ vccd1 _03112_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11819__A1 game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10089_ _04284_ _04296_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__nor2_1
X_14966_ game.CPU.walls.rand_wall.count_luck\[5\] game.CPU.walls.rand_wall.count_luck\[4\]
+ game.CPU.walls.rand_wall.count_luck\[1\] _08721_ _08727_ vssd1 vssd1 vccd1 vccd1
+ _08743_ sky130_fd_sc_hd__a311o_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16705_ net186 _02486_ net106 _02568_ net1533 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[147\]
+ sky130_fd_sc_hd__a32o_1
X_13917_ net862 game.CPU.applesa.ab.check_walls.above.walls\[157\] _03463_ net938
+ _07790_ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__a221o_1
XFILLER_0_199_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19216__CLK net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17685_ _03062_ _03068_ _03069_ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__nor3_1
X_14897_ net1105 _08414_ vssd1 vssd1 vccd1 vccd1 _08674_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_334_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19424_ clknet_leaf_39_clk game.writer.tracker.next_frame\[19\] net1330 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_348_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16636_ net156 _02535_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__nor2_1
X_13848_ game.writer.tracker.frame\[565\] net836 net671 game.writer.tracker.frame\[568\]
+ vssd1 vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__o22a_1
XANTENNA__16456__B _02328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_256_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19355_ clknet_leaf_71_clk game.CPU.applesa.twoapples.absxs.next_head\[0\] vssd1
+ vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.x_final\[0\] sky130_fd_sc_hd__dfxtp_1
X_16567_ net210 net150 _02415_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_26_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10785__A game.CPU.applesa.ab.absxs.body_y\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13779_ _07651_ _07652_ net496 vssd1 vssd1 vccd1 vccd1 _07653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_312_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Left_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18306_ net621 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
X_15518_ _01517_ _01539_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__and2_1
XANTENNA__19366__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19286_ clknet_leaf_68_clk net533 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.y_final\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16498_ game.writer.tracker.frame\[65\] _02433_ _02443_ net127 vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[65\] sky130_fd_sc_hd__a22o_1
XANTENNA__17183__A1 _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13419__S1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18237_ net649 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
X_15449_ _08917_ _01474_ _01475_ _08925_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__o22a_1
XANTENNA__16472__A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16930__A1 _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15733__A2 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13744__B2 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18168_ net632 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
XANTENNA__10558__A1 game.CPU.applesa.ab.absxs.body_x\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10558__B2 game.CPU.applesa.ab.absxs.body_x\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold403 game.writer.tracker.frame\[219\] vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_345_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17119_ net186 _02524_ net76 _02708_ net1999 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[421\]
+ sky130_fd_sc_hd__a32o_1
Xhold414 game.writer.tracker.frame\[334\] vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12952__C1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15088__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold425 game.writer.tracker.frame\[115\] vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold436 game.writer.tracker.frame\[357\] vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12505__A game.CPU.applesa.ab.absxs.body_x\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18099_ net639 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13100__S net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold447 game.writer.tracker.frame\[396\] vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_269_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold458 game.CPU.randy.f1.a1.count\[15\] vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 game.writer.tracker.frame\[3\] vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ net1115 net1116 _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_267_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_284_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12224__B net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout905 _03200_ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__buf_4
XFILLER_0_96_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17238__A2 _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_84_Left_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout916 net918 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_8
Xfanout927 net928 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__buf_2
XFILLER_0_244_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09872_ net1093 _03258_ _03324_ net1159 _04109_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__a221o_1
XANTENNA__10025__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout938 net940 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_8
Xfanout949 net950 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_8
XANTENNA__16997__A1 _02477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_224_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16997__B2 game.writer.tracker.frame\[336\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09533__B game.CPU.applesa.ab.check_walls.above.walls\[73\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16461__A3 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12240__A game.CPU.applesa.ab.check_walls.above.walls\[151\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_356_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12483__B2 game.CPU.applesa.ab.absxs.body_y\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_353_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout454_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19700__RESET_B net1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19709__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout242_X net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout621_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout719_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ net1093 game.CPU.applesa.ab.absxs.body_x\[54\] vssd1 vssd1 vccd1 vccd1 _03549_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_307_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09237_ game.CPU.applesa.ab.check_walls.above.walls\[196\] vssd1 vssd1 vccd1 vccd1
+ _03486_ sky130_fd_sc_hd__inv_2
XANTENNA__18733__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19859__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16921__A1 _02289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16382__A _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1151_X net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1249_X net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13735__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12538__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09168_ game.CPU.applesa.ab.check_walls.above.walls\[67\] vssd1 vssd1 vccd1 vccd1
+ _03417_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout990_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12943__C1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09099_ game.CPU.applesa.ab.absxs.body_y\[27\] vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__inv_2
XANTENNA__09708__B game.CPU.applesa.ab.absxs.body_y\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_309_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_287_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13010__S net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11130_ _03237_ net406 vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__xnor2_1
XANTENNA__18883__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12134__B net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14160__A1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13594__S0 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17229__A2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ _03280_ net323 vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14160__B2 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16437__B1 _02398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ net1163 game.CPU.applesa.out_random_2\[4\] vssd1 vssd1 vccd1 vccd1 _04220_
+ sky130_fd_sc_hd__nand2_2
XANTENNA__16988__A1 _02470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10721__A1 game.CPU.applesa.ab.absxs.body_y\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14820_ game.CPU.randy.counter1.count\[15\] _08624_ net139 vssd1 vssd1 vccd1 vccd1
+ _08627_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_327_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16452__A3 _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__B net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_240_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11277__A2 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14751_ game.CPU.randy.counter1.count1\[16\] game.CPU.randy.counter1.count1\[15\]
+ _08571_ vssd1 vssd1 vccd1 vccd1 _08575_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11963_ net814 net303 _05845_ _05849_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_263_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13702_ _07574_ _07575_ net487 vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__mux2_1
XANTENNA__19441__RESET_B net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10914_ _04383_ _04472_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__or2_1
X_17470_ _02897_ _02898_ _02893_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__a21o_1
XANTENNA__19389__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11894_ net821 net303 vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__or2_1
X_14682_ _08509_ _08519_ vssd1 vssd1 vccd1 vccd1 _08521_ sky130_fd_sc_hd__nor2_1
XANTENNA__14215__A2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16276__B net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16421_ _02248_ net235 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__or2_2
X_13633_ game.writer.tracker.frame\[49\] game.writer.tracker.frame\[51\] game.writer.tracker.frame\[52\]
+ game.writer.tracker.frame\[50\] net977 net1024 vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__mux4_1
X_10845_ _03505_ game.CPU.randy.counter1.count\[8\] _03504_ game.CPU.randy.counter1.count1\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_128_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19140_ net1187 _00182_ _00811_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[185\]
+ sky130_fd_sc_hd__dfrtp_2
X_16352_ net2043 net734 _02337_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[25\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_39_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17165__A1 _02458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13564_ net219 _07429_ _07434_ _07437_ net276 vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__o221a_1
X_10776_ game.CPU.applesa.ab.absxs.body_y\[64\] _04679_ _04680_ game.CPU.applesa.ab.absxs.body_y\[60\]
+ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10788__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16563__Y _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12309__B net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15303_ game.CPU.applesa.twomode.number\[6\] _08846_ vssd1 vssd1 vccd1 vccd1 _08851_
+ sky130_fd_sc_hd__or2_1
X_19071_ net1185 _00106_ _00742_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_12515_ _06382_ _06387_ _06390_ _06391_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__or4b_1
XFILLER_0_164_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13495_ _07054_ _07056_ _07066_ _07055_ net705 net497 vssd1 vssd1 vccd1 vccd1 _07369_
+ sky130_fd_sc_hd__mux4_1
X_16283_ net248 _02285_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__or2_2
XANTENNA__16912__A1 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_298_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13726__A1 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18022_ net663 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__inv_2
XANTENNA__12529__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17180__A4 _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15234_ game.CPU.applesa.normal1.number\[7\] _08794_ vssd1 vssd1 vccd1 vccd1 _08797_
+ sky130_fd_sc_hd__xor2_1
X_12446_ game.CPU.applesa.ab.absxs.body_y\[90\] net517 vssd1 vssd1 vccd1 vccd1 _06323_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_251_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12934__C1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_301_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_300_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ net1227 net1253 game.CPU.walls.rand_wall.x_final\[1\] vssd1 vssd1 vccd1 vccd1
+ _00199_ sky130_fd_sc_hd__and3_1
X_12377_ game.CPU.applesa.ab.absxs.body_x\[113\] net378 net520 game.CPU.applesa.ab.absxs.body_y\[114\]
+ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__o22a_1
XANTENNA__09618__B game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_288_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14116_ net984 net785 vssd1 vssd1 vccd1 vccd1 _07990_ sky130_fd_sc_hd__xor2_1
X_11328_ _05196_ _05211_ _05216_ _05208_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__or4b_2
X_19973_ clknet_leaf_41_clk game.writer.tracker.next_frame\[568\] net1331 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[568\] sky130_fd_sc_hd__dfrtp_1
X_15096_ net1205 net1232 game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1
+ vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__and3_1
XFILLER_0_293_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12044__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18924_ clknet_leaf_5_clk net4 _00608_ vssd1 vssd1 vccd1 vccd1 game.CPU.left_button.sync1.Q
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14151__A1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14047_ net1071 game.CPU.applesa.ab.check_walls.above.walls\[192\] vssd1 vssd1 vccd1
+ vccd1 _07921_ sky130_fd_sc_hd__xor2_1
X_11259_ game.CPU.applesa.ab.absxs.body_x\[39\] net545 net542 game.CPU.applesa.ab.absxs.body_y\[37\]
+ _05111_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__o221a_1
XFILLER_0_238_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18012__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09634__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18855_ clknet_leaf_0_clk _01246_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11883__B net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16979__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_340_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14273__A1_N net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12331__Y game.CPU.applesa.twoapples.absxs.next_head\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17806_ _01541_ _03141_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18606__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18786_ clknet_leaf_3_clk game.CPU.state1.Qn\[0\] _00523_ vssd1 vssd1 vccd1 vccd1
+ game.CPU.clock1.game_state\[0\] sky130_fd_sc_hd__dfstp_4
X_15998_ _03431_ net270 net341 _03433_ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a22o_1
XANTENNA__14454__A2 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17737_ game.CPU.applesa.ab.count\[2\] game.CPU.applesa.ab.count\[1\] _03099_ vssd1
+ vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__nand3_1
X_14949_ game.CPU.walls.rand_wall.count_luck\[3\] _08725_ vssd1 vssd1 vccd1 vccd1
+ _08726_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_341_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09330__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09330__B2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17668_ game.CPU.kyle.L1.cnt_500hz\[13\] _03056_ _03057_ vssd1 vssd1 vccd1 vccd1
+ _01259_ sky130_fd_sc_hd__o21a_1
XFILLER_0_323_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14206__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19407_ clknet_leaf_48_clk game.writer.tracker.next_frame\[2\] net1294 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16619_ net68 _02518_ _02526_ net1923 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[103\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_46_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15090__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18756__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17599_ _03009_ _03015_ net582 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19338_ clknet_leaf_72_clk _01354_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.count_luck\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13965__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13965__B2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17156__A1 _02436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_176_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_351_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12219__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11123__B net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19269_ clknet_leaf_7_clk _00057_ _00899_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_344_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16903__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09022_ game.CPU.applesa.ab.absxs.body_x\[51\] vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10962__B net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold200 game.writer.tracker.frame\[165\] vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 game.writer.tracker.frame\[291\] vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout202_A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09528__B game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12235__A game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold222 game.writer.tracker.frame\[234\] vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold233 game.writer.tracker.frame\[394\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 game.CPU.applesa.twoapples.y_final\[1\] vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 game.writer.tracker.frame\[181\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold266 game.writer.tracker.frame\[405\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold277 game.CPU.randy.counter1.count\[10\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold288 game.writer.tracker.frame\[168\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__B2 game.CPU.applesa.ab.absxs.body_y\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold299 game.writer.tracker.frame\[382\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13576__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout702 net707 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09924_ net1079 _04163_ _04164_ _04156_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__o31a_1
XFILLER_0_284_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout713 net714 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__buf_2
XANTENNA__14450__A game.CPU.applesa.ab.absxs.body_y\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout724 net725 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_187_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1111_A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout735 net738 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1209_A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout746 _04450_ vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_4
XANTENNA__19952__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20044_ game.wr vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11793__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_244_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09855_ net1131 game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1 _04098_
+ sky130_fd_sc_hd__nand2_1
Xfanout757 game.CPU.applesa.twomode.counter vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input7_A gpio_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout571_A net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 game.CPU.applesa.ab.apple_possible\[2\] vssd1 vssd1 vccd1 vccd1 net768
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_304_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout779 game.CPU.applesa.ab.apple_possible\[0\] vssd1 vssd1 vccd1 vccd1 net779
+ sky130_fd_sc_hd__buf_4
XANTENNA_fanout669_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09786_ net1097 game.CPU.applesa.ab.check_walls.above.walls\[145\] vssd1 vssd1 vccd1
+ vccd1 _04029_ sky130_fd_sc_hd__or2_1
XANTENNA__19531__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14445__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13102__C1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11259__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout836_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_X net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_65_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_3_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09321__A1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09321__B2 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_202_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19681__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_327_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10630_ net933 game.CPU.applesa.ab.absxs.body_x\[53\] vssd1 vssd1 vccd1 vccd1 _04683_
+ sky130_fd_sc_hd__and2_1
XANTENNA__13956__A1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13956__B2 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17147__A1 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12129__B net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11033__B net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10561_ game.CPU.applesa.ab.absxs.body_x\[20\] _04645_ _04652_ game.CPU.applesa.ab.absxs.body_x\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_153_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13169__C1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12300_ _06184_ _06185_ _06182_ _06183_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__a211o_1
XANTENNA__13708__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13280_ game.writer.tracker.frame\[462\] game.writer.tracker.frame\[463\] net1010
+ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__mux2_1
XANTENNA__09719__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10492_ _04614_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout993_X net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11719__B1 game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_310_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09388__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12231_ net815 net550 vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__and2_1
XFILLER_0_295_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09388__B2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12392__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_287_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12162_ _06046_ _06047_ _06048_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__or3b_2
XPHY_EDGE_ROW_269_Right_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_229_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19061__CLK net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ game.CPU.applesa.ab.absxs.body_y\[35\] net396 vssd1 vssd1 vccd1 vccd1 _05003_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__14998__C game.CPU.applesa.ab.check_walls.above.walls\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16970_ _02435_ net96 _02661_ net1839 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[319\]
+ sky130_fd_sc_hd__a22o_1
X_12093_ game.CPU.applesa.ab.check_walls.above.walls\[100\] net554 vssd1 vssd1 vccd1
+ vccd1 _05980_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_208_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18629__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11044_ _03265_ net319 vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__xnor2_1
X_15921_ game.CPU.applesa.ab.check_walls.above.walls\[131\] net457 vssd1 vssd1 vccd1
+ vccd1 _01933_ sky130_fd_sc_hd__nor2_1
XFILLER_0_263_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13319__S0 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18640_ clknet_leaf_59_clk _01057_ _00377_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[38\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16425__A3 _02390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09560__B2 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15852_ game.CPU.applesa.ab.absxs.body_y\[96\] net455 vssd1 vssd1 vccd1 vccd1 _01864_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__16558__Y _02486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14436__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14803_ game.CPU.randy.counter1.count\[9\] game.CPU.randy.counter1.count\[8\] _08612_
+ vssd1 vssd1 vccd1 vccd1 _08616_ sky130_fd_sc_hd__and3_1
XFILLER_0_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11208__B net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18571_ clknet_leaf_62_clk _00991_ _00308_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13644__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15783_ _03267_ net352 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__xnor2_1
X_12995_ game.writer.tracker.frame\[514\] game.writer.tracker.frame\[515\] net1008
+ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_258_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16287__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_56_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_188_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17522_ net1243 _02924_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__or2_1
XANTENNA__16718__C _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14734_ game.CPU.randy.counter1.count1\[10\] _08561_ vssd1 vssd1 vccd1 vccd1 _08564_
+ sky130_fd_sc_hd__or2_1
X_11946_ net798 net305 vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__xor2_1
XANTENNA__16189__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__A2 game.CPU.applesa.ab.absxs.body_y\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14519__B _08392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17453_ _02807_ _02881_ _02814_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__a21oi_1
X_14665_ _08487_ _04356_ _04347_ vssd1 vssd1 vccd1 vccd1 _08504_ sky130_fd_sc_hd__and3b_1
X_11877_ net747 _05235_ _05764_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11670__A2 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_253_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16404_ net240 net167 _02279_ _02284_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__and4_4
XANTENNA__11224__A game.CPU.applesa.ab.absxs.body_y\[38\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13616_ game.writer.tracker.frame\[317\] game.writer.tracker.frame\[319\] game.writer.tracker.frame\[320\]
+ game.writer.tracker.frame\[318\] net979 net1034 vssd1 vssd1 vccd1 vccd1 _07490_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17138__A1 _02405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10828_ game.CPU.walls.enable_in2 net1243 _04734_ vssd1 vssd1 vccd1 vccd1 _00011_
+ sky130_fd_sc_hd__mux2_1
X_17384_ _02812_ _02813_ _02777_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__a21oi_1
X_14596_ _08455_ net741 _08454_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[2\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_54_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12039__B net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_345_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19123_ net1183 _00163_ _00794_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[168\]
+ sky130_fd_sc_hd__dfrtp_4
X_16335_ net240 net236 _02325_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__or3_4
X_13547_ game.writer.tracker.frame\[77\] game.writer.tracker.frame\[79\] game.writer.tracker.frame\[80\]
+ game.writer.tracker.frame\[78\] net974 net999 vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__mux4_1
XFILLER_0_326_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_298_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10759_ game.CPU.applesa.ab.absxs.body_y\[97\] net263 _04719_ game.CPU.applesa.ab.absxs.body_y\[93\]
+ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__a22o_1
XANTENNA__18007__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16897__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19054_ net1192 _00286_ _00725_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[99\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09629__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16266_ _02271_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__inv_2
X_13478_ net508 _07351_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__or2_1
XANTENNA__12326__Y game.CPU.applesa.twoapples.absxs.next_head\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18005_ net613 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__inv_2
XFILLER_0_313_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15217_ game.CPU.applesa.normal1.number\[4\] _08778_ vssd1 vssd1 vccd1 vccd1 _08783_
+ sky130_fd_sc_hd__or2_1
XANTENNA__19404__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12429_ game.CPU.applesa.ab.absxs.body_x\[100\] net384 vssd1 vssd1 vccd1 vccd1 _06306_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09348__B game.CPU.applesa.ab.absxs.body_y\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_285_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16197_ _02029_ _02030_ _02032_ _02033_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__or4_1
XANTENNA__16649__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_301_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15148_ net1210 net1236 game.CPU.applesa.ab.check_walls.above.walls\[176\] vssd1
+ vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__and3_1
XANTENNA__17310__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_236_Right_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_291_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_264_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19956_ clknet_leaf_43_clk game.writer.tracker.next_frame\[551\] net1305 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[551\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14270__A game.CPU.applesa.ab.absxs.body_y\[50\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15079_ net1211 net1237 game.CPU.applesa.ab.check_walls.above.walls\[107\] vssd1
+ vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__and3_1
XANTENNA__19554__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_206_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15085__B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18907_ clknet_leaf_9_clk _01274_ _00591_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_19887_ clknet_leaf_27_clk game.writer.tracker.next_frame\[482\] net1311 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[482\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12502__B net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17074__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__B2 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ net1126 net788 vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__nand2_1
X_18838_ clknet_leaf_0_clk _01229_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16468__Y _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09571_ net919 game.CPU.applesa.ab.absxs.body_x\[78\] game.CPU.applesa.ab.absxs.body_y\[79\]
+ net906 _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__a221o_1
XANTENNA__11118__B net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18769_ clknet_leaf_50_clk _01186_ _00506_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[71\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13635__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12438__B2 game.CPU.applesa.ab.absxs.body_y\[106\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_47_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_353_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09811__B game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17377__A1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10957__B net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14429__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout152_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11661__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10464__A3 _04594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11134__A game.CPU.applesa.ab.absxs.body_y\[69\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17129__A1 net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_217_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16644__B _02404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10973__A game.CPU.applesa.ab.absxs.body_y\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_A net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1061_A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1159_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09005_ game.CPU.applesa.ab.absxs.body_x\[105\] vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14363__A1 game.CPU.applesa.ab.absxs.body_x\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_277_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13879__A2_N game.CPU.applesa.ab.check_walls.above.walls\[106\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14363__B2 game.CPU.applesa.ab.absxs.body_y\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout205_X net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1326_A net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_306_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_203_Right_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout510 net511 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13323__C1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout521 net522 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_2
Xfanout532 _06212_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_4
X_09907_ net1100 _04147_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__or2_1
Xfanout543 _04815_ vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout953_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout554 net555 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_4
Xfanout565 _04461_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_4
XANTENNA__17065__B1 _02689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__A1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18921__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout576 _08937_ vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_2
XANTENNA__09542__B2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__A game.CPU.applesa.ab.check_walls.above.walls\[67\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_20027_ net1277 vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
X_09838_ net1093 _03253_ game.CPU.applesa.ab.absxs.body_y\[107\] net908 _04080_ vssd1
+ vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__o221a_1
Xfanout587 net591 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__buf_2
Xfanout598 net625 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__buf_2
XFILLER_0_308_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16812__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11028__B net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15723__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12839__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14179__X _08053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ net1129 net802 vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__16538__C _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16114__A2_N game.CPU.applesa.ab.absxs.body_y\[69\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11800_ game.CPU.applesa.ab.check_walls.above.walls\[198\] net304 _05682_ _05686_
+ _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12443__A2_N net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10500__X _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12780_ game.writer.tracker.frame\[96\] game.writer.tracker.frame\[97\] net1012 vssd1
+ vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__mux2_2
XFILLER_0_96_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_317_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11731_ net800 net311 vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14450_ game.CPU.applesa.ab.absxs.body_y\[12\] net994 vssd1 vssd1 vccd1 vccd1 _08324_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11662_ game.CPU.applesa.ab.check_walls.above.walls\[123\] net761 vssd1 vssd1 vccd1
+ vccd1 _05551_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_354_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_338_Right_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13401_ _06866_ _06879_ net685 vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__mux2_1
XANTENNA__19427__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11979__A game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10613_ net1080 _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__nor2_2
X_14381_ game.CPU.applesa.ab.absxs.body_y\[81\] net861 net856 game.CPU.applesa.ab.absxs.body_y\[83\]
+ _08250_ vssd1 vssd1 vccd1 vccd1 _08255_ sky130_fd_sc_hd__o221a_1
X_11593_ game.CPU.applesa.ab.check_walls.above.walls\[104\] net775 vssd1 vssd1 vccd1
+ vccd1 _05482_ sky130_fd_sc_hd__xor2_1
XFILLER_0_354_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_289_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16120_ game.CPU.applesa.ab.check_walls.above.walls\[177\] net475 net347 _03476_
+ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__a2bb2o_1
X_13332_ net480 _06924_ _07205_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10544_ game.CPU.applesa.ab.absxs.body_x\[36\] _04642_ _04643_ game.CPU.applesa.ab.absxs.body_x\[32\]
+ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__a22o_1
XANTENNA__10612__B1 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16051_ game.CPU.applesa.ab.absxs.body_x\[100\] net273 vssd1 vssd1 vccd1 vccd1 _02063_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_161_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13788__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13263_ net477 _07136_ net681 vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__a21o_1
X_10475_ _03263_ _04601_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__nor2_1
XFILLER_0_269_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12365__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19577__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15002_ net1223 net1251 game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1
+ vccd1 vccd1 _00219_ sky130_fd_sc_hd__and3_1
XANTENNA__19874__RESET_B net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13562__C1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12214_ game.CPU.applesa.ab.check_walls.above.walls\[175\] net424 vssd1 vssd1 vccd1
+ vccd1 _06100_ sky130_fd_sc_hd__nor2_1
X_13194_ game.writer.tracker.frame\[402\] game.writer.tracker.frame\[403\] net1039
+ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19810_ clknet_leaf_39_clk game.writer.tracker.next_frame\[405\] net1353 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[405\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09781__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ game.CPU.applesa.ab.check_walls.above.walls\[190\] net289 net295 net781 vssd1
+ vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09781__B2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12162__X _06049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_263_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14090__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13314__C1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10300__A_N game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16953_ _02404_ net95 _02657_ net1737 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[306\]
+ sky130_fd_sc_hd__a22o_1
X_19741_ clknet_leaf_25_clk game.writer.tracker.next_frame\[336\] net1320 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[336\] sky130_fd_sc_hd__dfrtp_2
X_12076_ _05958_ _05959_ _05960_ _05962_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__or4_1
XANTENNA__12668__A1 net1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ _03264_ net326 vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__xnor2_1
X_15904_ _01907_ _01909_ _01914_ _01915_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__or4_1
X_19672_ clknet_leaf_32_clk game.writer.tracker.next_frame\[267\] net1285 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[267\] sky130_fd_sc_hd__dfrtp_1
X_16884_ _02272_ net119 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__nand2_4
XFILLER_0_218_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11340__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14409__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18623_ clknet_leaf_11_clk _01040_ _00360_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[105\]
+ sky130_fd_sc_hd__dfrtp_4
X_15835_ game.CPU.applesa.ab.absxs.body_y\[108\] net452 vssd1 vssd1 vccd1 vccd1 _01847_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15192__Y _00016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_204_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13712__S0 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18554_ clknet_leaf_45_clk _00977_ net1300 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.cmd_num\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13093__A1 game.writer.tracker.frame\[241\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15766_ _01772_ _01773_ _01775_ _01777_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__or4_1
XFILLER_0_63_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12978_ net702 _06617_ _06614_ net210 vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__o211a_1
XANTENNA__14249__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11037__A2_N net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17505_ net1264 _02933_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__nor2_1
X_14717_ _08551_ _08552_ net54 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__and3b_1
X_11929_ game.CPU.applesa.ab.check_walls.above.walls\[189\] net306 net300 game.CPU.applesa.ab.check_walls.above.walls\[190\]
+ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18485_ net638 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__inv_2
X_15697_ game.CPU.applesa.ab.absxs.body_x\[31\] net457 net438 game.CPU.applesa.ab.absxs.body_y\[30\]
+ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__a22o_1
XFILLER_0_170_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17436_ game.CPU.modea.Qa\[0\] _02845_ _02850_ _02859_ vssd1 vssd1 vccd1 vccd1 _02866_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14648_ _04350_ _04555_ _08486_ vssd1 vssd1 vccd1 vccd1 _08487_ sky130_fd_sc_hd__nor3_1
XFILLER_0_184_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_345_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_333_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _05781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_305_Right_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18733__Q game.CPU.applesa.ab.absxs.body_x\[115\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_39 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17367_ _02796_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__inv_2
X_14579_ game.CPU.clock1.counter\[9\] game.CPU.clock1.counter\[14\] game.CPU.clock1.counter\[16\]
+ _03520_ vssd1 vssd1 vccd1 vccd1 _08441_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10793__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19106_ net1180 _00145_ _00777_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[151\]
+ sky130_fd_sc_hd__dfrtp_2
X_16318_ net1965 net722 _02312_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[16\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__10603__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09359__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17298_ net1968 net723 _02756_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[552\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_259_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19037_ net1193 _00268_ _00708_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[82\]
+ sky130_fd_sc_hd__dfrtp_4
X_16249_ net186 net171 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__nand2_4
XFILLER_0_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_212_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15808__B net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10906__A1 game.CPU.applesa.enable_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16098__A1 game.CPU.applesa.ab.absxs.body_x\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09772__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16098__B2 game.CPU.applesa.ab.absxs.body_y\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13609__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09772__B2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19939_ clknet_leaf_38_clk game.writer.tracker.next_frame\[534\] net1331 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[534\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16479__X _02429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_345_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_301_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18200__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09822__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ _03859_ _03860_ _03865_ _03858_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__a211o_1
XFILLER_0_207_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18908__Q game.CPU.applesa.ab.absxs.body_y\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_223_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout367_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13344__A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13703__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ net1141 game.CPU.applesa.ab.absxs.body_y\[62\] vssd1 vssd1 vccd1 vccd1 _03797_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_179_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_328_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18556__SET_B net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09485_ net920 game.CPU.applesa.ab.check_walls.above.walls\[186\] _03481_ net1157
+ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout155_X net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout534_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18643__Q game.CPU.applesa.ab.absxs.body_y\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1064_X net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_312_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12595__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_305_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11311__B net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_249_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16390__A _02252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1329_X net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12347__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10260_ game.CPU.applesa.ab.XMAX\[1\] _04441_ net746 net774 game.CPU.applesa.ab.XMAX\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__o32a_1
XFILLER_0_239_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_284_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10191_ net1097 _04383_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_7_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_226_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1305 net1306 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__clkbuf_2
Xfanout1316 net1323 vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__clkbuf_4
Xfanout1327 net1334 vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__buf_2
XFILLER_0_319_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1338 net1341 vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 game.CPU.walls.rand_wall.abduyd.next_wall\[5\] vssd1 vssd1 vccd1 vccd1
+ net340 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12142__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1349 net1351 vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_255_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17038__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout351 net352 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_148_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout362 net363 vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_323_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout373 net374 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_2
X_13950_ net881 game.CPU.applesa.ab.check_walls.above.walls\[129\] _03449_ net983
+ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__o22a_1
Xfanout384 net385 vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__buf_4
XANTENNA_fanout68_X net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 _05604_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12901_ game.writer.tracker.frame\[20\] game.writer.tracker.frame\[21\] net1024 vssd1
+ vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__mux2_1
XANTENNA__09732__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13881_ _07750_ _07752_ _07754_ vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__and3_1
XFILLER_0_213_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10878__A game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13254__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15620_ game.CPU.applesa.ab.check_walls.above.walls\[87\] net433 vssd1 vssd1 vccd1
+ vccd1 _01632_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_335_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12832_ game.writer.tracker.frame\[282\] game.writer.tracker.frame\[283\] net1017
+ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__mux2_1
XANTENNA__16800__A3 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_295_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _01497_ _01537_ _08936_ _01491_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a211o_1
XFILLER_0_201_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12763_ _06634_ _06583_ _06587_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__and3b_1
XFILLER_0_271_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_237_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14502_ _08373_ _08374_ _08375_ _08372_ vssd1 vssd1 vccd1 vccd1 _08376_ sky130_fd_sc_hd__a211o_1
X_11714_ net811 net311 vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__nand2_1
X_18270_ net649 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
X_15482_ _08903_ _08918_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__or2_2
XANTENNA__18817__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12694_ _06565_ _06567_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__and2_1
XANTENNA__14024__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16284__B _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17221_ net67 net142 net119 _02736_ net1553 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[495\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_204_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19298__D net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14433_ _08304_ _08305_ _08306_ vssd1 vssd1 vccd1 vccd1 _08307_ sky130_fd_sc_hd__or3_1
XFILLER_0_126_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_343_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11645_ _05488_ _05504_ _05520_ _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__and4_1
XFILLER_0_154_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17152_ _02429_ net58 _02717_ net1772 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[445\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_342_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14364_ game.CPU.applesa.ab.absxs.body_x\[103\] net873 net962 _03294_ _08233_ vssd1
+ vssd1 vccd1 vccd1 _08238_ sky130_fd_sc_hd__a221o_1
XFILLER_0_330_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11576_ game.CPU.applesa.ab.check_walls.above.walls\[134\] net254 vssd1 vssd1 vccd1
+ vccd1 _05465_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_5_clk_X clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16103_ _03354_ net454 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__nand2_1
X_13315_ net240 _07182_ _07187_ _07188_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__a31o_1
XANTENNA__11221__B net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17083_ net206 _02386_ net57 _02697_ net1832 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[396\]
+ sky130_fd_sc_hd__a32o_1
X_10527_ game.CPU.applesa.ab.absxs.body_x\[55\] _04609_ _04637_ game.CPU.applesa.ab.absxs.body_x\[51\]
+ vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__a22o_1
XANTENNA__16867__A3 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14295_ _03240_ net1050 net864 game.CPU.applesa.ab.absxs.body_y\[53\] vssd1 vssd1
+ vccd1 vccd1 _08169_ sky130_fd_sc_hd__a22o_1
X_16034_ game.CPU.applesa.ab.absxs.body_x\[45\] net474 vssd1 vssd1 vccd1 vccd1 _02046_
+ sky130_fd_sc_hd__and2_1
X_13246_ _07116_ _07117_ _07118_ _07119_ net487 net682 vssd1 vssd1 vccd1 vccd1 _07120_
+ sky130_fd_sc_hd__mux4_1
X_10458_ _04580_ _04592_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__or2_2
XANTENNA__09907__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15628__B net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_248_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13177_ game.writer.tracker.frame\[442\] game.writer.tracker.frame\[443\] net1040
+ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_296_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10389_ net919 game.CPU.apple_location\[2\] game.CPU.apple_location\[3\] net925 vssd1
+ vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12333__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_261_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12128_ net832 net555 vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__or2_1
XANTENNA__17292__A3 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17985_ net628 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__inv_2
XANTENNA__16299__X _02299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19724_ clknet_leaf_35_clk game.writer.tracker.next_frame\[319\] net1346 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[319\] sky130_fd_sc_hd__dfrtp_1
X_16936_ _02369_ net92 _02652_ net1490 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[294\]
+ sky130_fd_sc_hd__a22o_1
X_12059_ game.CPU.applesa.ab.check_walls.above.walls\[197\] net387 vssd1 vssd1 vccd1
+ vccd1 _05946_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15644__A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18020__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16459__B net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09642__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19655_ clknet_leaf_22_clk game.writer.tracker.next_frame\[250\] net1343 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[250\] sky130_fd_sc_hd__dfrtp_1
X_16867_ net152 _02422_ net107 _02628_ net1671 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[249\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__16252__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18606_ clknet_leaf_69_clk _01023_ _00343_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[88\]
+ sky130_fd_sc_hd__dfrtp_4
X_15818_ game.CPU.applesa.ab.absxs.body_x\[90\] net465 vssd1 vssd1 vccd1 vccd1 _01830_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_337_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19586_ clknet_leaf_36_clk game.writer.tracker.next_frame\[181\] net1351 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[181\] sky130_fd_sc_hd__dfrtp_1
X_16798_ _02478_ net103 _02600_ net1763 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[208\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14263__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18537_ net611 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__inv_2
X_15749_ game.CPU.applesa.ab.check_walls.above.walls\[2\] net468 vssd1 vssd1 vccd1
+ vccd1 _01761_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_259_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10824__A0 net1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09270_ game.CPU.applesa.enable_in vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__inv_2
X_18468_ net652 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19742__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17419_ _02841_ _02848_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__and2_1
X_18399_ net617 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12508__A game.CPU.applesa.ab.absxs.body_y\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13103__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12577__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11412__A game.CPU.applesa.ab.check_walls.above.walls\[115\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17504__A1 game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12041__A2 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload54_A clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11131__B net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19892__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12942__S net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_259_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout115_A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_348_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12329__B1 net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_259_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10970__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14442__B net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11823__D_N _05710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17268__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09745__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09745__B2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1024_A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13829__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ game.CPU.applesa.ab.absxs.body_x\[84\] vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_299_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout484_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09552__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19272__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A _08799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16243__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_A _04442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ net1093 game.CPU.applesa.ab.absxs.body_x\[118\] vssd1 vssd1 vccd1 vccd1 _03849_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_197_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16794__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11068__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__B _05194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ net901 net813 game.CPU.applesa.ab.check_walls.above.walls\[75\] net928 vssd1
+ vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_167_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout537_X net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout916_A net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1279_X net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09468_ net1091 _03229_ _03297_ net1146 _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__a221o_1
XFILLER_0_241_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_325_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12418__A game.CPU.applesa.ab.absxs.body_x\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09399_ net1130 game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1 vccd1
+ vccd1 _03642_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11322__A game.CPU.applesa.ab.check_walls.above.walls\[68\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11430_ game.CPU.applesa.ab.check_walls.above.walls\[27\] net763 vssd1 vssd1 vccd1
+ vccd1 _05319_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_151_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10043__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11361_ game.CPU.applesa.ab.check_walls.above.walls\[39\] net261 vssd1 vssd1 vccd1
+ vccd1 _05250_ sky130_fd_sc_hd__xor2_1
XANTENNA__13780__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16849__A3 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_232_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Left_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13100_ _06935_ _06937_ net687 vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__mux2_1
X_10312_ game.CPU.randy.f1.a1.count\[12\] game.CPU.randy.f1.a1.count\[11\] game.CPU.randy.f1.a1.count\[10\]
+ _04494_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__and4_1
XANTENNA__15448__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11292_ _05063_ _05070_ _05175_ _05181_ _05105_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__o311a_1
X_14080_ net963 game.CPU.applesa.ab.check_walls.above.walls\[93\] vssd1 vssd1 vccd1
+ vccd1 _07954_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14352__B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09736__A1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13031_ net698 _06875_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__or2_1
X_10243_ _03213_ game.CPU.luck1.Qa\[0\] _04435_ net846 vssd1 vssd1 vccd1 vccd1 _04436_
+ sky130_fd_sc_hd__o31a_1
XANTENNA__13532__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09736__B2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12153__A game.CPU.applesa.ab.check_walls.above.walls\[135\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ net1168 game.CPU.applesa.ab.apple_possible\[5\] vssd1 vssd1 vccd1 vccd1 _04367_
+ sky130_fd_sc_hd__nand2_2
Xfanout1102 net1104 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__buf_4
XANTENNA__17274__A3 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1113 game.CPU.applesa.ab.snake_head_x\[0\] vssd1 vssd1 vccd1 vccd1 net1113
+ sky130_fd_sc_hd__buf_4
Xfanout1124 game.CPU.bodymain1.main.score\[0\] vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__clkbuf_4
XANTENNA__19615__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1135 net1138 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__buf_4
XANTENNA__11992__A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17770_ game.CPU.applesa.twoapples.count_luck\[6\] _03121_ _03109_ vssd1 vssd1 vccd1
+ vccd1 _01355_ sky130_fd_sc_hd__o21a_1
Xfanout1146 net1152 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__buf_4
X_14982_ net1224 net1250 game.CPU.applesa.ab.check_walls.above.walls\[10\] vssd1 vssd1
+ vccd1 vccd1 _00187_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_89_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1157 game.CPU.applesa.ab.snake_head_y\[0\] vssd1 vssd1 vccd1 vccd1 net1157
+ sky130_fd_sc_hd__clkbuf_8
Xfanout170 _02255_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_218_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14493__B1 _08164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1168 net1169 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16279__B _08400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1179 net1190 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__buf_2
X_16721_ _02257_ _02427_ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__nor2_1
XANTENNA__09462__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13933_ net873 game.CPU.applesa.ab.check_walls.above.walls\[35\] _03399_ net986 vssd1
+ vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__a22o_1
XANTENNA__13391__S1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11846__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19440_ clknet_leaf_43_clk game.writer.tracker.next_frame\[35\] net1303 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[35\] sky130_fd_sc_hd__dfrtp_1
X_16652_ net168 net155 net69 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__and3_2
X_13864_ net281 _07732_ _07737_ net485 vssd1 vssd1 vccd1 vccd1 _07738_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16785__A2 _02460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19765__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_241_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15603_ game.CPU.applesa.ab.check_walls.above.walls\[113\] net471 net346 _03440_
+ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__a2bb2o_1
X_12815_ _06687_ _06688_ net501 vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_215_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19371_ clknet_leaf_71_clk _01377_ _00952_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location2\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11216__B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16583_ net1759 _02500_ _02502_ net126 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[91\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15911__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13795_ game.writer.tracker.frame\[391\] net711 net838 game.writer.tracker.frame\[389\]
+ vssd1 vssd1 vccd1 vccd1 _07669_ sky130_fd_sc_hd__o22a_1
X_18322_ net615 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_303_Left_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15534_ _01523_ _01546_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__nor2_1
X_12746_ game.writer.tracker.frame\[80\] game.writer.tracker.frame\[81\] net999 vssd1
+ vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__mux2_2
XFILLER_0_96_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_316_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18253_ net644 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
X_15465_ _08936_ _01491_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__nor2_1
X_12677_ net879 net875 vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__nor2_2
XFILLER_0_56_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12328__A net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17204_ net156 _02365_ net71 net715 vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__o31a_1
XANTENNA__11232__A game.CPU.applesa.ab.absxs.body_x\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12559__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14416_ _08284_ _08289_ vssd1 vssd1 vccd1 vccd1 _08290_ sky130_fd_sc_hd__or2_1
X_11628_ net566 _05508_ _05511_ _05513_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__a211o_1
X_18184_ net609 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_170_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13220__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15396_ game.writer.updater.commands.cmd_num\[1\] game.writer.updater.commands.cmd_num\[3\]
+ game.writer.updater.commands.cmd_num\[4\] game.writer.updater.commands.cmd_num\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08938_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_303_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_122_Left_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17135_ net165 _02396_ _02690_ _02713_ game.writer.tracker.frame\[432\] vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.next_frame\[432\] sky130_fd_sc_hd__a32o_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13771__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14347_ game.CPU.applesa.ab.absxs.body_y\[33\] net960 vssd1 vssd1 vccd1 vccd1 _08221_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12615__X _06492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11559_ game.CPU.applesa.ab.check_walls.above.walls\[196\] net251 vssd1 vssd1 vccd1
+ vccd1 _05448_ sky130_fd_sc_hd__xnor2_1
XANTENNA__18015__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 game.writer.tracker.frame\[131\] vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10585__A2 _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19145__CLK net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold618 game.writer.tracker.frame\[353\] vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13508__C1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold629 game.writer.tracker.frame\[328\] vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
X_17066_ _02241_ _02634_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__nor2_2
X_14278_ _08146_ _08151_ vssd1 vssd1 vccd1 vccd1 _08152_ sky130_fd_sc_hd__or2_1
XANTENNA__16170__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_312_Left_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09727__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16017_ game.CPU.applesa.ab.absxs.body_x\[38\] net469 vssd1 vssd1 vccd1 vccd1 _02029_
+ sky130_fd_sc_hd__xnor2_1
X_13229_ _07086_ _07102_ net247 vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__a21o_1
XANTENNA__13523__A2 _07391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19295__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16473__B2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17968_ net668 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_181_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13287__B2 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_131_Left_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14484__B1 _08357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09372__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19707_ clknet_leaf_32_clk game.writer.tracker.next_frame\[302\] net1284 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[302\] sky130_fd_sc_hd__dfrtp_1
X_16919_ _02342_ _02643_ net559 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17899_ net657 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__inv_2
XANTENNA__12510__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19638_ clknet_leaf_28_clk game.writer.tracker.next_frame\[233\] net1287 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[233\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16776__A2 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_321_Left_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_342_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11126__B net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19569_ clknet_leaf_32_clk game.writer.tracker.next_frame\[164\] net1296 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[164\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09322_ _03556_ _03557_ _03559_ _03560_ _03564_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_319_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10965__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10273__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_307_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09253_ game.CPU.randy.counter1.count\[12\] vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__inv_2
XANTENNA__10273__B2 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09184_ game.CPU.applesa.ab.check_walls.above.walls\[100\] vssd1 vssd1 vccd1 vccd1
+ _03433_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13211__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12014__A2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16652__B net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09966__A1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10981__A game.CPU.applesa.ab.absxs.body_x\[73\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1141_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout118_X net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1239_A net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09547__A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14172__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19638__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout699_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10045__X _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_281_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17256__A3 _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16464__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12701__A _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ game.CPU.kyle.L1.nextState\[3\] vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_145_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14475__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18662__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19788__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_320_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_230_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10930_ _03357_ net535 vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16767__A2 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_316_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_205_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_252_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15731__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ _03500_ game.CPU.randy.counter1.count1\[13\] game.CPU.randy.counter1.count1\[12\]
+ _03501_ _04757_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ game.CPU.applesa.ab.absxs.body_x\[109\] net378 net372 game.CPU.applesa.ab.absxs.body_x\[110\]
+ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_84_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_292_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ net276 _07445_ net238 vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_26_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10792_ net937 game.CPU.applesa.ab.absxs.body_y\[44\] net562 _04727_ vssd1 vssd1
+ vccd1 vccd1 _01003_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_234_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14347__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12531_ game.CPU.applesa.ab.absxs.body_x\[97\] net376 net369 _03325_ _06407_ vssd1
+ vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__o221a_1
XANTENNA__17939__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17192__A2 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19168__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15250_ net264 vssd1 vssd1 vccd1 vccd1 _08811_ sky130_fd_sc_hd__inv_2
X_12462_ game.CPU.applesa.ab.absxs.body_y\[110\] net520 vssd1 vssd1 vccd1 vccd1 _06339_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_23_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_340_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14201_ game.CPU.applesa.ab.absxs.body_x\[64\] net888 net985 _03336_ vssd1 vssd1
+ vccd1 vccd1 _08075_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11413_ game.CPU.applesa.ab.check_walls.above.walls\[114\] net767 vssd1 vssd1 vccd1
+ vccd1 _05302_ sky130_fd_sc_hd__xor2_2
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15181_ game.CPU.bodymain1.main.score\[4\] _04577_ _08756_ net1115 vssd1 vssd1 vccd1
+ vccd1 _08757_ sky130_fd_sc_hd__o31ai_1
X_12393_ game.CPU.applesa.ab.absxs.body_y\[25\] net527 net517 game.CPU.applesa.ab.absxs.body_y\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__a22o_1
XANTENNA__10567__A2 _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14132_ net987 game.CPU.applesa.ab.check_walls.above.walls\[44\] vssd1 vssd1 vccd1
+ vccd1 _08006_ sky130_fd_sc_hd__xor2_1
XANTENNA__16152__B1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344_ net808 net258 _05232_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_293_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13505__A2 _07375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14063_ net1071 _03456_ _03457_ net1052 _07930_ vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__a221o_1
X_18940_ net1176 _00079_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number_out\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_277_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11275_ net1270 net399 net412 game.CPU.applesa.ab.absxs.body_x\[61\] vssd1 vssd1
+ vccd1 vccd1 _05165_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11516__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13014_ game.writer.tracker.frame\[532\] game.writer.tracker.frame\[533\] net1021
+ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_265_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_245_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10226_ game.CPU.applesa.ab.count_luck\[6\] game.CPU.applesa.ab.count_luck\[7\] vssd1
+ vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__or2_1
XANTENNA__15906__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18871_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[1\] _00566_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19662__Q game.writer.tracker.frame\[257\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16455__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17822_ _03147_ _03148_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__nand2_1
XANTENNA__10830__S _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ _03220_ _04349_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_167_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_233_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14466__B1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 game.CPU.start_pause_button1.eD1.D vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09192__A game.CPU.applesa.ab.check_walls.above.walls\[115\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17753_ _03110_ _03111_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__nor2_1
X_14965_ _03488_ game.CPU.luck1.Qa\[0\] _08741_ _04253_ vssd1 vssd1 vccd1 vccd1 _08742_
+ sky130_fd_sc_hd__o31a_1
X_10088_ _04214_ _04222_ _04294_ _04292_ _04288_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__o32a_1
XANTENNA__11819__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__A game.CPU.applesa.ab.absxs.body_x\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16704_ _02322_ _02561_ net735 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__o21a_1
X_13916_ net1062 game.CPU.applesa.ab.check_walls.above.walls\[153\] vssd1 vssd1 vccd1
+ vccd1 _07790_ sky130_fd_sc_hd__xor2_1
XANTENNA__15922__A game.CPU.applesa.ab.check_walls.above.walls\[135\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17684_ game.CPU.walls.rand_wall.count_luck\[3\] _03066_ vssd1 vssd1 vccd1 vccd1
+ _03069_ sky130_fd_sc_hd__nor2_1
XFILLER_0_226_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14896_ _08670_ _08672_ vssd1 vssd1 vccd1 vccd1 _08673_ sky130_fd_sc_hd__nor2_1
XFILLER_0_202_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_334_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19423_ clknet_leaf_39_clk game.writer.tracker.next_frame\[18\] net1330 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[18\] sky130_fd_sc_hd__dfrtp_1
X_16635_ net172 _02479_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__or2_4
XFILLER_0_186_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13847_ game.writer.tracker.frame\[569\] game.writer.tracker.frame\[571\] game.writer.tracker.frame\[572\]
+ game.writer.tracker.frame\[570\] net982 net1022 vssd1 vssd1 vccd1 vccd1 _07721_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__15641__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13442__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16566_ net216 _02415_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__and2_2
X_19354_ clknet_leaf_71_clk _01364_ _00939_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.logic_enable
+ sky130_fd_sc_hd__dfstp_1
X_13778_ game.writer.tracker.frame\[145\] game.writer.tracker.frame\[147\] game.writer.tracker.frame\[148\]
+ game.writer.tracker.frame\[146\] net977 net1023 vssd1 vssd1 vccd1 vccd1 _07652_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_256_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12875__S0 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__B _04630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15517_ _08039_ _01514_ _01471_ _08028_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__a211o_1
X_18305_ net641 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
X_12729_ game.writer.tracker.frame\[102\] game.writer.tracker.frame\[103\] net995
+ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19285_ clknet_leaf_69_clk game.CPU.applesa.ab.good_spot_next vssd1 vssd1 vccd1 vccd1
+ game.CPU.applesa.ab.good_spot sky130_fd_sc_hd__dfxtp_1
X_16497_ net158 _02438_ _02442_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__a21o_1
XANTENNA__17183__A2 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18236_ net650 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
XFILLER_0_217_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15448_ net943 net954 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__nand2_1
XFILLER_0_331_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14544__Y _08416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16472__B net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19837__Q game.writer.tracker.frame\[432\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16930__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18741__Q game.CPU.applesa.ab.absxs.body_x\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11897__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18167_ net628 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15379_ _08900_ _08915_ vssd1 vssd1 vccd1 vccd1 _08921_ sky130_fd_sc_hd__or2_1
XANTENNA__11755__A1 game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17118_ net186 _02521_ net81 _02708_ net2017 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[420\]
+ sky130_fd_sc_hd__a32o_1
Xhold404 game.writer.tracker.frame\[491\] vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15800__A1_N game.CPU.applesa.ab.absxs.body_y\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09367__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_345_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold415 game.writer.tracker.frame\[68\] vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15088__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18098_ net611 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__inv_2
XANTENNA__16143__B1 net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold426 game.writer.tracker.frame\[308\] vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold437 game.writer.tracker.frame\[216\] vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12505__B net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold448 game.writer.tracker.frame\[198\] vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16694__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold459 game.writer.tracker.frame\[374\] vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
X_17049_ _02415_ _02678_ _02685_ net1844 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[374\]
+ sky130_fd_sc_hd__a22o_1
X_09940_ _04175_ _04177_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__nor2_1
XFILLER_0_269_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14560__X _08427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_267_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18685__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout906 net907 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__buf_4
XFILLER_0_110_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_337_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17238__A3 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19930__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09871_ net1132 game.CPU.applesa.ab.absxs.body_y\[111\] vssd1 vssd1 vccd1 vccd1 _04114_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_209_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout917 net918 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15816__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_244_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout928 _03192_ vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_4
XFILLER_0_284_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout939 net940 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkload17_A clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16446__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_209_Left_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16997__A2 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_224_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16487__X _02435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_252_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13680__A1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09884__B1 _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_356_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1091_A game.CPU.applesa.ab.snake_head_x\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10976__A game.CPU.applesa.ab.absxs.body_y\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_278_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout447_A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1189_A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13432__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14167__B net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09305_ net1111 game.CPU.applesa.ab.absxs.body_x\[52\] vssd1 vssd1 vccd1 vccd1 _03548_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16663__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_218_Left_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout614_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17174__A2 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10797__A2 _04690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_334_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_302_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09236_ game.CPU.applesa.ab.check_walls.above.walls\[194\] vssd1 vssd1 vccd1 vccd1
+ _03485_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_334_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_30_clk_X clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_334_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16921__A2 _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16382__B _02359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13498__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_302_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19460__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09167_ net816 vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13291__S0 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_X net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16134__B1 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ game.CPU.applesa.ab.absxs.body_y\[32\] vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_309_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout983_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12415__B net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16685__A1 _02267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_45_clk_X clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12104__A2_N net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout95_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11060_ game.CPU.applesa.ab.absxs.body_y\[27\] net396 vssd1 vssd1 vccd1 vccd1 _04950_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__17229__A3 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14160__A2 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_227_Left_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15726__B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16437__A1 game.writer.tracker.frame\[49\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10011_ net897 _04218_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16437__B2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09283__Y _03528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14448__B1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16988__A2 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15661__A2_N net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10721__A2 _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11318__Y _05207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_327_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_231_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15742__A game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750_ _08573_ _08574_ net55 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_240_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ game.CPU.applesa.ab.check_walls.above.walls\[68\] net394 net309 net815 vssd1
+ vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09875__B1 _04019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13701_ game.writer.tracker.frame\[465\] game.writer.tracker.frame\[467\] game.writer.tracker.frame\[468\]
+ game.writer.tracker.frame\[466\] net974 net1011 vssd1 vssd1 vccd1 vccd1 _07575_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09740__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913_ net416 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.next_head\[0\] sky130_fd_sc_hd__inv_2
XANTENNA__19828__RESET_B net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14681_ _08506_ _08508_ vssd1 vssd1 vccd1 vccd1 _08520_ sky130_fd_sc_hd__or2_1
X_11893_ _05777_ _05778_ _05780_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__and3_1
XANTENNA__14358__A game.CPU.applesa.ab.absxs.body_y\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16420_ net115 net164 net53 _02384_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[44\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_345_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_343_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13632_ game.writer.tracker.frame\[55\] net712 net675 game.writer.tracker.frame\[56\]
+ _07505_ vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__o221a_1
XANTENNA__16276__C _02280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10844_ _03507_ game.CPU.randy.counter1.count1\[6\] _03509_ game.CPU.randy.counter1.count1\[5\]
+ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_236_Left_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16351_ net1993 net734 _02337_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[24\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_183_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18558__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13563_ net500 _07430_ _07431_ net201 vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10775_ game.CPU.applesa.ab.absxs.body_y\[65\] _04679_ _04680_ game.CPU.applesa.ab.absxs.body_y\[61\]
+ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__a22o_1
XANTENNA__19803__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15302_ game.CPU.applesa.twomode.number\[2\] _08844_ vssd1 vssd1 vccd1 vccd1 _08850_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__10788__A2 game.CPU.applesa.ab.absxs.body_y\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_212_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19070_ net1185 _00105_ _00741_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[115\]
+ sky130_fd_sc_hd__dfrtp_4
X_12514_ game.CPU.applesa.ab.absxs.body_x\[75\] net531 net519 game.CPU.applesa.ab.absxs.body_y\[74\]
+ _06385_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__o221a_1
X_16282_ _02279_ _02284_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13494_ _07049_ _07050_ _07060_ _07051_ net706 net497 vssd1 vssd1 vccd1 vccd1 _07368_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_217_Right_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18021_ net663 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15233_ _00019_ _08793_ _08794_ _08795_ _08796_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__o32a_1
XANTENNA__18561__Q game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12445_ _06321_ _06317_ _06316_ _06319_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__and4b_1
XFILLER_0_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_251_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11510__A game.CPU.applesa.ab.check_walls.above.walls\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12934__B1 _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14524__C _07742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15164_ net1225 net1252 game.CPU.walls.rand_wall.x_final\[0\] vssd1 vssd1 vccd1 vccd1
+ _00088_ sky130_fd_sc_hd__and3_1
XANTENNA__16125__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19953__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ game.CPU.applesa.ab.absxs.body_x\[112\] net383 vssd1 vssd1 vccd1 vccd1 _06253_
+ sky130_fd_sc_hd__and2_1
XANTENNA__16676__A1 game.writer.tracker.frame\[129\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15476__X net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14115_ net1069 game.CPU.applesa.ab.check_walls.above.walls\[168\] vssd1 vssd1 vccd1
+ vccd1 _07989_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11327_ net814 net257 _05214_ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__a211o_1
X_19972_ clknet_leaf_41_clk game.writer.tracker.next_frame\[567\] net1331 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[567\] sky130_fd_sc_hd__dfrtp_1
X_15095_ net1203 net1229 game.CPU.applesa.ab.check_walls.above.walls\[123\] vssd1
+ vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__and3_1
XANTENNA__14240__A2_N net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ net949 game.CPU.applesa.ab.check_walls.above.walls\[198\] vssd1 vssd1 vccd1
+ vccd1 _07920_ sky130_fd_sc_hd__xor2_1
XANTENNA__09915__A game.CPU.applesa.clk_body vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18923_ clknet_leaf_4_clk net1407 _00607_ vssd1 vssd1 vccd1 vccd1 game.CPU.left_button.eD1.Q2
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14151__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15636__B net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11258_ _05085_ _05086_ _05087_ _05091_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19392__Q game.CPU.bad_collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10209_ _04398_ _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__xor2_1
XFILLER_0_207_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15629__A2_N net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12341__A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18854_ clknet_leaf_6_clk _01245_ _00564_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09634__B game.CPU.applesa.ab.absxs.body_y\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11189_ _05073_ _05074_ _05075_ _05076_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__a22o_1
XANTENNA__16979__A2 _02454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_340_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_234_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17805_ net943 net954 _06573_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__and3_1
XANTENNA__12060__B net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18785_ clknet_leaf_10_clk _01202_ _00522_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_15997_ game.CPU.applesa.ab.check_walls.above.walls\[100\] net451 net439 net803 vssd1
+ vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a22o_1
XANTENNA__13111__A0 game.writer.tracker.frame\[144\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15652__A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17736_ _03099_ _03100_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__nor2_1
X_14948_ game.CPU.walls.rand_wall.count_luck\[1\] game.CPU.walls.rand_wall.count_luck\[0\]
+ game.CPU.walls.rand_wall.count_luck\[2\] vssd1 vssd1 vccd1 vccd1 _08725_ sky130_fd_sc_hd__a21o_1
XFILLER_0_167_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19333__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16467__B _02376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09650__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19569__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10476__B2 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17667_ game.CPU.kyle.L1.cnt_500hz\[13\] _03056_ net194 vssd1 vssd1 vccd1 vccd1 _03057_
+ sky130_fd_sc_hd__a21boi_1
X_14879_ game.CPU.walls.abc.number\[3\] game.CPU.walls.abc.number\[7\] game.CPU.walls.abc.counter
+ vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__mux2_1
XANTENNA__16600__A1 _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_334_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19406_ clknet_leaf_47_clk game.writer.tracker.next_frame\[1\] net1294 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[1\] sky130_fd_sc_hd__dfrtp_1
X_16618_ net145 net124 _02369_ _02526_ net1868 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[102\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__13414__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17598_ game.CPU.kyle.L1.cnt_20ms\[4\] _03002_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16549_ net196 _02314_ _02316_ net240 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__o22a_4
XANTENNA__19483__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19337_ clknet_leaf_72_clk _01353_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.count_luck\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13965__A2 game.CPU.applesa.ab.check_walls.above.walls\[177\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17156__A2 net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_351_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13900__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09649__X _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19268_ clknet_leaf_7_clk _00056_ _00898_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13178__A0 _07048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17561__C1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16903__A2 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09021_ game.CPU.applesa.ab.absxs.body_x\[59\] vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ net666 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__inv_2
XANTENNA__14914__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19199_ clknet_leaf_67_clk _01308_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_331_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11420__A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09097__A game.CPU.applesa.ab.absxs.body_y\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold201 game.writer.tracker.frame\[399\] vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14390__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold212 game.writer.tracker.frame\[283\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 game.writer.tracker.frame\[508\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12235__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16667__B2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold234 game.writer.tracker.frame\[94\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 game.writer.tracker.frame\[270\] vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 game.writer.tracker.frame\[196\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold267 game.writer.tracker.frame\[404\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18203__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 game.writer.tracker.frame\[235\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09825__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09923_ net922 net1262 vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__nor2_1
Xfanout703 net707 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__buf_2
Xhold289 game.writer.tracker.frame\[472\] vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout714 net726 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_113_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14450__B net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_272_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout725 net726 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_187_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout397_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout736 net737 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_4
X_20043_ net1367 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout747 net748 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_2
X_09854_ _04088_ _04089_ _04090_ _04096_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__or4_2
Xfanout758 game.CPU.applesa.normal1.counter vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1104_A game.CPU.applesa.ab.snake_head_x\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_304_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10703__A2 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17092__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09785_ net1097 game.CPU.applesa.ab.check_walls.above.walls\[145\] vssd1 vssd1 vccd1
+ vccd1 _04028_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout185_X net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout564_A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19992__RESET_B net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_319_Right_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_339_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_72_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19921__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18646__Q game.CPU.applesa.ab.absxs.body_y\[52\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18700__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19826__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1094_X net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11154__X _05044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16198__A3 _02208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_313_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1359_X net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10560_ game.CPU.applesa.ab.absxs.body_x\[21\] _04645_ _04652_ game.CPU.applesa.ab.absxs.body_x\[17\]
+ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__a22o_1
XANTENNA__18850__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19976__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09219_ game.CPU.applesa.ab.check_walls.above.walls\[165\] vssd1 vssd1 vccd1 vccd1
+ _03468_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10645__S _04690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10491_ _04580_ _04583_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__nand2_2
XANTENNA__12426__A game.CPU.applesa.ab.absxs.body_y\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11719__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ net815 net550 vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__or2_1
XANTENNA__14381__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16107__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_295_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout986_X net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19206__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_287_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12161_ game.CPU.applesa.ab.check_walls.above.walls\[39\] net296 net291 net822 vssd1
+ vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout98_X net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11112_ _03275_ net319 vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_248_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11984__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12092_ net804 net388 vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11043_ game.CPU.applesa.ab.absxs.body_x\[81\] net414 vssd1 vssd1 vccd1 vccd1 _04933_
+ sky130_fd_sc_hd__xnor2_1
X_15920_ game.CPU.applesa.ab.check_walls.above.walls\[131\] net457 vssd1 vssd1 vccd1
+ vccd1 _01932_ sky130_fd_sc_hd__and2_1
XFILLER_0_290_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19356__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17083__A1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13319__S1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11048__Y _04938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15851_ game.CPU.applesa.ab.absxs.body_x\[98\] net466 vssd1 vssd1 vccd1 vccd1 _01863_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_164_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_290_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15472__A _01454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14802_ _08614_ _08615_ vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15782_ game.CPU.applesa.ab.absxs.body_y\[75\] net433 vssd1 vssd1 vccd1 vccd1 _01794_
+ sky130_fd_sc_hd__xnor2_1
X_18570_ clknet_leaf_8_clk _00990_ _00307_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_12994_ game.writer.tracker.frame\[566\] game.writer.tracker.frame\[567\] net1021
+ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09848__B1 game.CPU.applesa.ab.absxs.body_y\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17521_ _02825_ net426 _02840_ _02878_ _02823_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__a311o_1
X_14733_ game.CPU.randy.counter1.count1\[10\] _08561_ vssd1 vssd1 vccd1 vccd1 _08563_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_244_Left_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11945_ net799 net390 vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17452_ _02787_ _02801_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__nor2_1
XFILLER_0_184_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14664_ game.CPU.randy.counter1.count1\[9\] _08500_ _08502_ game.CPU.randy.counter1.count1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _08503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11876_ net747 _05235_ _05236_ net569 vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_129_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16574__Y _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16403_ net1752 _02371_ _02374_ net135 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[39\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13615_ game.writer.tracker.frame\[313\] game.writer.tracker.frame\[315\] game.writer.tracker.frame\[316\]
+ game.writer.tracker.frame\[314\] net979 net1034 vssd1 vssd1 vccd1 vccd1 _07489_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_253_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11999__X _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10827_ game.CPU.walls.enable_in2 game.CPU.modea.Qa\[0\] _04735_ vssd1 vssd1 vccd1
+ vccd1 _00008_ sky130_fd_sc_hd__mux2_1
X_17383_ net1114 net1115 game.CPU.bodymain1.main.score\[7\] vssd1 vssd1 vccd1 vccd1
+ _02813_ sky130_fd_sc_hd__o21a_1
XANTENNA__11224__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14595_ game.CPU.clock1.counter\[1\] game.CPU.clock1.counter\[0\] game.CPU.clock1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _08455_ sky130_fd_sc_hd__and3_1
XANTENNA__17138__A2 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11958__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16334_ _02245_ _02284_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__nand2_1
X_19122_ net1182 _00162_ _00793_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[167\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13546_ _07417_ _07418_ _07419_ net278 net241 vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10758_ game.CPU.applesa.ab.absxs.body_y\[98\] net263 _04719_ game.CPU.applesa.ab.absxs.body_y\[94\]
+ vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_299_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16897__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19053_ net1192 _00285_ _00724_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[98\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16265_ net173 net159 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__nand2_4
X_13477_ _07130_ _07155_ net700 vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__mux2_1
XANTENNA__11252__A2_N net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09629__B game.CPU.applesa.ab.absxs.body_x\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10689_ game.CPU.applesa.ab.absxs.body_y\[100\] _04595_ _04708_ game.CPU.applesa.ab.absxs.body_y\[96\]
+ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15216_ _08782_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__inv_2
X_18004_ net634 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__inv_2
X_12428_ net1265 net531 vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_341_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_253_Left_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14372__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16196_ _01628_ _01629_ _02207_ _01625_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__a211o_1
XFILLER_0_112_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16649__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13580__B1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15147_ net1214 net1239 game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1
+ vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__and3_1
X_12359_ game.CPU.applesa.ab.absxs.body_y\[46\] net520 vssd1 vssd1 vccd1 vccd1 _06236_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18023__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14551__A net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17310__A2 _02535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11894__B net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19955_ clknet_leaf_43_clk game.writer.tracker.next_frame\[550\] net1303 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[550\] sky130_fd_sc_hd__dfrtp_1
X_15078_ net1211 net1237 game.CPU.applesa.ab.check_walls.above.walls\[106\] vssd1
+ vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_264_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14270__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13167__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_284_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_206_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14029_ net959 _03468_ net787 net852 vssd1 vssd1 vccd1 vccd1 _07903_ sky130_fd_sc_hd__a22o_1
X_18906_ clknet_leaf_9_clk _01273_ _00590_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_254_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19886_ clknet_leaf_27_clk game.writer.tracker.next_frame\[481\] net1311 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[481\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15085__C game.CPU.applesa.ab.check_walls.above.walls\[113\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17074__A1 _02456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18837_ clknet_leaf_0_clk _01228_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__19849__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09570_ net919 game.CPU.applesa.ab.absxs.body_x\[78\] game.CPU.applesa.ab.absxs.body_x\[77\]
+ net914 vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_262_Left_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12438__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18768_ clknet_leaf_53_clk _01185_ _00505_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[70\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17719_ game.CPU.applesa.ab.count_luck\[1\] _03086_ net1535 vssd1 vssd1 vccd1 vccd1
+ _03090_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_353_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18699_ clknet_leaf_60_clk _01116_ _00436_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17801__S net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__A game.CPU.applesa.ab.check_walls.above.walls\[113\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18873__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19999__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16484__Y _02432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_275_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11835__A2_N net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11134__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12945__S net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_217_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17129__A2 _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13494__S0 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout145_A net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11949__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13630__A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10973__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_271_Left_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12246__A game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout312_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_A game.CPU.applesa.x\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ game.CPU.applesa.ab.absxs.body_x\[106\] vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__inv_2
XANTENNA__14363__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_277_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout100_X net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1221_A game.CPU.walls.rand_wall.start_enable vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_306_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1319_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09801__A1_N net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09555__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout681_A _06600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout500 net503 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14180__B net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 net515 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_228_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout779_A game.CPU.applesa.ab.apple_possible\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09906_ net1100 _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__nand2_1
Xfanout522 _06214_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__buf_2
Xfanout533 net537 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_4
XFILLER_0_272_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_245_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1107_X net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_4
XANTENNA__17065__A1 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout555 _04777_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_4
Xfanout566 _04460_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_4
XANTENNA__10688__A1 game.CPU.applesa.ab.absxs.body_y\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_20026_ net1277 vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
X_09837_ net908 game.CPU.applesa.ab.absxs.body_y\[107\] game.CPU.applesa.ab.absxs.body_y\[104\]
+ net893 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__o2bb2a_1
Xfanout577 net578 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09542__A2 game.CPU.applesa.ab.XMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout588 net590 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_4
XANTENNA__11309__B net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_A game.CPU.applesa.y\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout599 net625 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout567_X net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ net1129 net802 vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_197_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout58_A net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09290__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_240_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09699_ net1086 game.CPU.applesa.ab.check_walls.above.walls\[59\] vssd1 vssd1 vccd1
+ vccd1 _03942_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_317_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13016__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11325__A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11730_ net801 net301 vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__nand2_1
XFILLER_0_324_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_354_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_260_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11044__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11661_ game.CPU.applesa.ab.check_walls.above.walls\[12\] net252 _05544_ _05545_
+ _05546_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__o2111a_1
XANTENNA__14051__A1 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14051__B2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13400_ _07272_ _07273_ net484 vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10612_ _04591_ _04615_ _04625_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__a21o_4
XANTENNA__11979__B net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14380_ game.CPU.applesa.ab.absxs.body_x\[80\] net886 net852 game.CPU.applesa.ab.absxs.body_y\[82\]
+ _08253_ vssd1 vssd1 vccd1 vccd1 _08254_ sky130_fd_sc_hd__o221a_1
XFILLER_0_153_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11592_ net775 _05480_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_289_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13331_ net500 _06735_ net695 vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__a21o_1
X_10543_ game.CPU.applesa.ab.absxs.body_x\[37\] _04642_ _04643_ game.CPU.applesa.ab.absxs.body_x\[33\]
+ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__a22o_1
XANTENNA__17947__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12156__A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16050_ game.CPU.applesa.ab.absxs.body_y\[100\] net454 vssd1 vssd1 vccd1 vccd1 _02062_
+ sky130_fd_sc_hd__xnor2_1
X_13262_ game.writer.tracker.frame\[484\] game.writer.tracker.frame\[485\] net1010
+ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__mux2_1
XANTENNA__14354__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10474_ _04603_ game.CPU.applesa.ab.absxs.body_x\[94\] _04601_ vssd1 vssd1 vccd1
+ vccd1 _01197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_269_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12365__A1 game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15001_ net1223 net1251 game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1
+ vccd1 vccd1 _00218_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_328_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12365__B2 game.CPU.applesa.ab.absxs.body_y\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12213_ _03474_ net421 vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ game.writer.tracker.frame\[404\] game.writer.tracker.frame\[405\] net1040
+ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12144_ _06028_ _06029_ _06030_ _06027_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__a211o_1
XANTENNA__09465__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14090__B game.CPU.applesa.ab.check_walls.above.walls\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_291_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12603__B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_263_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11059__X _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19740_ clknet_leaf_18_clk game.writer.tracker.next_frame\[335\] net1289 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[335\] sky130_fd_sc_hd__dfrtp_1
X_16952_ _02405_ _02638_ net729 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__o21a_1
XFILLER_0_285_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12075_ _05223_ _05225_ _05226_ _05227_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__or4_1
XANTENNA__13865__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11913__A1_N net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17056__A1 _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11026_ _03326_ net541 vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__nand2_1
X_15903_ _01906_ _01908_ _01910_ _01913_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__or4_1
X_19671_ clknet_leaf_32_clk game.writer.tracker.next_frame\[266\] net1292 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[266\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15914__B net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11219__B net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16883_ _02271_ _02634_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__nor2_1
XANTENNA__16298__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10123__B game.CPU.applesa.ab.good_collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_244_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13715__A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18622_ clknet_leaf_16_clk _01039_ _00359_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[104\]
+ sky130_fd_sc_hd__dfrtp_4
X_15834_ game.CPU.applesa.ab.absxs.body_x\[108\] net272 vssd1 vssd1 vccd1 vccd1 _01846_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09912__B net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18553_ clknet_leaf_45_clk _00976_ net1279 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.cmd_num\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_12977_ net213 _06648_ _06850_ net283 vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__a211o_1
X_15765_ _03285_ net344 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_231_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11235__A game.CPU.applesa.ab.absxs.body_x\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15930__A game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17504_ game.CPU.clock1.game_state\[0\] _02837_ _02822_ vssd1 vssd1 vccd1 vccd1 _02933_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11928_ net572 _05508_ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14716_ game.CPU.randy.counter1.count1\[4\] _08548_ vssd1 vssd1 vccd1 vccd1 _08552_
+ sky130_fd_sc_hd__or2_1
X_15696_ game.CPU.applesa.ab.absxs.body_y\[28\] net449 vssd1 vssd1 vccd1 vccd1 _01708_
+ sky130_fd_sc_hd__xnor2_1
X_18484_ net638 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__inv_2
XFILLER_0_234_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17435_ _02819_ _02823_ _02846_ _02855_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__or4_1
X_14647_ game.CPU.randy.f1.state\[4\] game.CPU.randy.f1.state\[5\] vssd1 vssd1 vccd1
+ vccd1 _08486_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11859_ net573 _05489_ _05495_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_318_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18018__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12053__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_29 _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ game.CPU.speed1.Qa\[2\] _08439_ _08438_ _08437_ _08436_ vssd1 vssd1 vccd1
+ vccd1 _08440_ sky130_fd_sc_hd__a2111o_1
X_17366_ net1117 _02795_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__or2_1
XANTENNA__10793__B _04690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12337__Y game.CPU.applesa.twoapples.absxs.next_head\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_19105_ net1181 _00144_ _00776_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[150\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13529_ game.writer.tracker.frame\[89\] game.writer.tracker.frame\[91\] game.writer.tracker.frame\[92\]
+ game.writer.tracker.frame\[90\] net979 net1018 vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__mux4_1
X_16317_ net1891 net722 _02312_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[15\]
+ sky130_fd_sc_hd__and3_1
X_17297_ net130 _02370_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12066__A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09600__A2_N game.CPU.applesa.ab.absxs.body_x\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16248_ net191 net169 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__nor2_1
X_19036_ net1192 _00267_ _00707_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[81\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__19521__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15542__A1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14345__A2 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_212_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13596__S net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16179_ _01759_ _01762_ _01764_ _01767_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__or4_1
XANTENNA__10367__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16098__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09375__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15096__B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19671__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19938_ clknet_leaf_42_clk game.writer.tracker.next_frame\[533\] net1326 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[533\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_254_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13856__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12659__A2 game.CPU.applesa.twoapples.absxs.next_head\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17047__A1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_184_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_345_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_242_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11129__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19869_ clknet_leaf_20_clk game.writer.tracker.next_frame\[464\] net1308 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[464\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_126_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_301_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09622_ net1160 _03379_ _03381_ net1131 _03864_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__a221o_1
XANTENNA__09822__B game.CPU.applesa.ab.absxs.body_x\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10968__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_223_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13344__B _06762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _03788_ _03789_ _03790_ _03795_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__or4_1
XANTENNA__16495__X _02441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout262_A _05195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11145__A game.CPU.applesa.ab.absxs.body_y\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_194_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09484_ _03724_ _03726_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_159_Left_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_336_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14456__A game.CPU.applesa.ab.absxs.body_x\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout148_X net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1171_A game.CPU.applesa.ab.YMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1269_A game.CPU.applesa.ab.absxs.body_x\[49\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18619__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_336_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13241__C1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_351_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_312_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_349_Left_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_310_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15558__Y net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16390__B net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18769__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13544__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14191__A game.CPU.applesa.ab.absxs.body_y\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1224_X net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_168_Left_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17286__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_284_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10190_ net1168 net769 vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_264_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1306 net1307 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__clkbuf_4
Xfanout1317 net1323 vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__clkbuf_4
Xfanout1328 net1329 vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__clkbuf_4
Xfanout330 _04647_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_2
Xfanout1339 net1341 vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17038__A1 _02238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout341 net342 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_8
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_6
XANTENNA__11727__A2_N net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_358_Left_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_255_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout363 _06218_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_323_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout374 _06210_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_6
Xfanout385 _06208_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_4
XANTENNA_fanout949_X net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12900_ game.writer.tracker.frame\[24\] game.writer.tracker.frame\[25\] net1025 vssd1
+ vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__mux2_1
Xfanout396 net400 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_4
XANTENNA__13535__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20009_ net1378 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
X_13880_ net880 game.CPU.applesa.ab.check_walls.above.walls\[106\] game.CPU.applesa.ab.check_walls.above.walls\[108\]
+ net867 _07753_ vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__o221a_1
XANTENNA__09732__B game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10530__B1 _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12831_ game.writer.tracker.frame\[284\] game.writer.tracker.frame\[285\] net1017
+ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_335_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_177_Left_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15550_ net576 _01455_ _01464_ _01538_ _01570_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__a311o_2
X_12762_ _06583_ _06587_ _06635_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_87_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_295_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_328_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17210__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ game.CPU.apple_location\[2\] net1053 vssd1 vssd1 vccd1 vccd1 _08375_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_237_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11713_ net811 net311 vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__or2_1
X_15481_ _08914_ _08921_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12693_ _06559_ _06560_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__xor2_4
XFILLER_0_204_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14024__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14024__B2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_351_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17220_ _02536_ net75 net557 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a21oi_1
X_14432_ _03281_ net1070 net869 game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1
+ vccd1 vccd1 _08306_ sky130_fd_sc_hd__a22o_1
XFILLER_0_166_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_355_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11644_ _05521_ _05530_ _05531_ _05532_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_159_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19544__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16852__Y _02623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17151_ _02428_ net58 _02717_ net1791 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[444\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_13_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14363_ game.CPU.applesa.ab.absxs.body_x\[102\] net878 net864 game.CPU.applesa.ab.absxs.body_y\[101\]
+ _08235_ vssd1 vssd1 vccd1 vccd1 _08237_ sky130_fd_sc_hd__a221o_1
X_11575_ game.CPU.applesa.ab.check_walls.above.walls\[134\] net254 vssd1 vssd1 vccd1
+ vccd1 _05464_ sky130_fd_sc_hd__or2_1
XANTENNA__17513__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16102_ game.CPU.applesa.ab.absxs.body_y\[16\] net341 vssd1 vssd1 vccd1 vccd1 _02114_
+ sky130_fd_sc_hd__nand2_1
X_13314_ _07167_ _07168_ _07172_ _07174_ net247 vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__o221a_2
XFILLER_0_220_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17082_ _02303_ _02693_ net725 vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__o21a_1
XFILLER_0_181_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10526_ net754 _04608_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__nor2_4
X_14294_ game.CPU.applesa.ab.absxs.body_x\[52\] net889 net994 _03308_ _08167_ vssd1
+ vssd1 vccd1 vccd1 _08168_ sky130_fd_sc_hd__a221o_1
XFILLER_0_220_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_186_Left_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16033_ game.CPU.applesa.ab.absxs.body_x\[45\] net474 vssd1 vssd1 vccd1 vccd1 _02045_
+ sky130_fd_sc_hd__nor2_1
X_13245_ game.writer.tracker.frame\[498\] game.writer.tracker.frame\[499\] net1016
+ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__mux2_1
XANTENNA__19694__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10457_ net1117 _03198_ _04358_ _04579_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__or4_2
XANTENNA__09195__A game.CPU.applesa.ab.check_walls.above.walls\[121\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ game.writer.tracker.frame\[446\] game.writer.tracker.frame\[447\] net1038
+ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_248_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10388_ net897 game.CPU.apple_location\[5\] _04538_ _04539_ net1263 vssd1 vssd1 vccd1
+ vccd1 _04540_ sky130_fd_sc_hd__o221a_1
XFILLER_0_236_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_261_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12127_ net832 net555 vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__nand2_1
X_17984_ net606 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
XANTENNA__17029__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19723_ clknet_leaf_35_clk game.writer.tracker.next_frame\[318\] net1346 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[318\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09923__A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16935_ _02370_ _02636_ net713 vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__o21a_1
X_12058_ _03486_ net555 vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15644__B net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16459__C _02415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ game.CPU.applesa.ab.absxs.body_y\[54\] net540 vssd1 vssd1 vccd1 vccd1 _04899_
+ sky130_fd_sc_hd__nor2_1
X_19654_ clknet_leaf_22_clk game.writer.tracker.next_frame\[249\] net1343 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[249\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09642__B game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16866_ _02545_ net99 net730 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__o21a_1
XANTENNA__16788__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16252__A2 _02252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_195_Left_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18605_ clknet_leaf_3_clk _00007_ _00342_ vssd1 vssd1 vccd1 vccd1 game.CPU.luck1.Qa\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_15817_ game.CPU.applesa.ab.absxs.body_y\[89\] net444 vssd1 vssd1 vccd1 vccd1 _01829_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__19074__CLK net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_337_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19585_ clknet_leaf_35_clk game.writer.tracker.next_frame\[180\] net1339 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[180\] sky130_fd_sc_hd__dfrtp_1
X_16797_ _02476_ net103 _02600_ net1573 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[207\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_245_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14263__A1 game.CPU.applesa.ab.absxs.body_x\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13697__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14263__B2 game.CPU.applesa.ab.absxs.body_x\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_181_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_247_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18536_ net628 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
X_15748_ game.CPU.applesa.ab.check_walls.above.walls\[2\] net468 vssd1 vssd1 vccd1
+ vccd1 _01760_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_259_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17201__A1 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10824__A1 net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18467_ net661 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_272_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15679_ _03385_ net334 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_261_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17418_ _02826_ _02847_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_334_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16960__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18398_ net617 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12508__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13774__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11412__B net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17349_ _03218_ net1259 vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__nand2_2
XANTENNA__18911__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16491__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14563__X _08429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14318__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_314_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15819__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_348_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload47_A clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19019_ net1196 _00248_ _00690_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[64\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_286_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout108_A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17268__A1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_239_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12243__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14117__A1_N game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08984_ game.CPU.applesa.ab.absxs.body_x\[85\] vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_299_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_270_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19417__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09552__B game.CPU.applesa.ab.absxs.body_x\[115\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16779__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ net1142 game.CPU.applesa.ab.absxs.body_y\[118\] vssd1 vssd1 vccd1 vccd1 _03848_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_155_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout644_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16666__A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09536_ net928 game.CPU.applesa.ab.check_walls.above.walls\[75\] net813 net901 vssd1
+ vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__19567__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16385__B net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ net1107 game.CPU.applesa.ab.absxs.body_x\[92\] vssd1 vssd1 vccd1 vccd1 _03710_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__14006__A1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout909_A _03199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1174_X net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14006__B2 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09398_ net1148 net806 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12418__B net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13765__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18591__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11322__B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09433__A1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09433__B2 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11360_ _05244_ _05245_ _05246_ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_10_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15729__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_277_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10311_ game.CPU.randy.f1.a1.count\[13\] game.CPU.randy.f1.a1.count\[9\] _04491_
+ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11291_ _04948_ _04949_ _05180_ _04894_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_325_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13030_ _06873_ _06888_ net698 vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__mux2_1
XANTENNA__17259__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ _04428_ _04434_ _04423_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_277_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12740__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10173_ _04364_ _04365_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1103 net1104 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__buf_4
XANTENNA_fanout80_X net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1114 game.CPU.bodymain1.main.score\[6\] vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_2
Xfanout1125 net1126 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__buf_4
XFILLER_0_218_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09743__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1136 net1138 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__buf_4
XANTENNA__11992__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1152 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__clkbuf_4
Xfanout160 _02256_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_206_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14981_ net1225 net1252 game.CPU.applesa.ab.check_walls.above.walls\[9\] vssd1 vssd1
+ vccd1 vccd1 _00176_ sky130_fd_sc_hd__and3_1
Xfanout1158 net1161 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__buf_4
Xfanout171 net172 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_245_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1169 game.CPU.applesa.ab.enable vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__clkbuf_2
X_16720_ _02343_ net99 net735 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__o21a_1
XFILLER_0_245_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout182 _03146_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
XANTENNA__09462__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13932_ _07802_ _07803_ _07804_ _07805_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__a22o_1
XANTENNA__17431__A1 net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16651_ _02415_ _02518_ _02543_ net1859 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[118\]
+ sky130_fd_sc_hd__a22o_1
X_13863_ game.writer.tracker.frame\[551\] net708 net671 game.writer.tracker.frame\[552\]
+ _07736_ vssd1 vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_18_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16785__A3 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12814_ _06684_ _06685_ net678 vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__mux2_1
X_15602_ _01610_ _01611_ _01612_ _01613_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__or4_1
X_19370_ clknet_leaf_71_clk _01376_ _00951_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13794_ net230 _07663_ _07667_ net286 vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__o211a_1
X_16582_ net195 _02297_ _02439_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18321_ net615 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__inv_2
X_12745_ _06569_ _06577_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__xnor2_1
X_15533_ _06562_ _01551_ _01505_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10806__B2 game.CPU.applesa.ab.absxs.body_y\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18934__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14096__A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11072__X _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11513__A game.CPU.applesa.ab.check_walls.above.walls\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_316_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15464_ _01464_ _01490_ _01487_ _01489_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__and4bb_1
X_18252_ net644 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
X_12676_ net883 _06549_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__or2_1
XFILLER_0_328_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17203_ net66 net122 net121 _02731_ net1517 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[482\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_231_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14415_ _08285_ _08286_ _08287_ _08288_ vssd1 vssd1 vccd1 vccd1 _08289_ sky130_fd_sc_hd__or4_1
XANTENNA__11232__B net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11627_ game.CPU.applesa.ab.check_walls.above.walls\[188\] net250 _05509_ net564
+ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__a221o_1
X_15395_ _03363_ game.writer.updater.commands.mode\[0\] vssd1 vssd1 vccd1 vccd1 _08937_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09424__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18183_ net610 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__inv_2
XANTENNA__09424__B2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17498__A1 game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17134_ _02394_ net72 net725 vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__o21a_1
X_14346_ _08217_ _08218_ _08219_ vssd1 vssd1 vccd1 vccd1 _08220_ sky130_fd_sc_hd__or3_1
X_11558_ net566 _05440_ _05446_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15639__B net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold608 game.writer.tracker.frame\[24\] vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11782__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17065_ net187 _02449_ _02689_ net1961 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[386\]
+ sky130_fd_sc_hd__a22o_1
X_10509_ game.CPU.applesa.ab.absxs.body_x\[70\] _04625_ _04626_ game.CPU.applesa.ab.absxs.body_x\[66\]
+ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__a22o_1
Xhold619 game.writer.tracker.frame\[100\] vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ _08148_ _08150_ vssd1 vssd1 vccd1 vccd1 _08151_ sky130_fd_sc_hd__nand2_1
XANTENNA__16170__A1 game.CPU.applesa.ab.absxs.body_x\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11489_ _05314_ _05331_ _05346_ _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__or4_1
XANTENNA__13603__S0 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire180_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16016_ net784 net451 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__xnor2_1
X_13228_ net215 _07101_ _07094_ net285 vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__a211o_1
XANTENNA__14181__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15655__A game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13159_ game.writer.tracker.frame\[154\] game.writer.tracker.frame\[155\] net1036
+ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18031__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_236_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09653__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_224_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18739__Q game.CPU.applesa.ab.absxs.body_x\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17967_ net668 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__inv_2
XFILLER_0_264_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_181_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_326_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_236_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19706_ clknet_leaf_31_clk game.writer.tracker.next_frame\[301\] net1284 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[301\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_224_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16918_ _02498_ net95 _02647_ net1881 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[281\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09372__B game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15093__C game.CPU.applesa.ab.check_walls.above.walls\[121\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17898_ net657 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19637_ clknet_leaf_28_clk game.writer.tracker.next_frame\[232\] net1287 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[232\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11407__B net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16849_ net131 _02391_ net122 _02620_ net1583 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[238\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_205_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_251_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_220_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13903__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19568_ clknet_leaf_48_clk game.writer.tracker.next_frame\[163\] net1296 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[163\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09321_ net1150 _03335_ _03336_ net1160 _03563_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__a221o_1
X_18519_ net581 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__inv_2
X_19499_ clknet_leaf_26_clk game.writer.tracker.next_frame\[94\] net1319 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[94\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09252_ game.CPU.randy.counter1.count\[13\] vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__inv_2
XANTENNA__11470__A1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16492__Y _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_192_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11142__B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09183_ game.CPU.applesa.ab.check_walls.above.walls\[99\] vssd1 vssd1 vccd1 vccd1
+ _03432_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout225_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16652__C net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09828__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09966__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10981__B net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09547__B game.CPU.applesa.ab.absxs.body_y\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12254__A net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1134_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_281_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1301_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10733__B1 _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16464__A2 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ game.CPU.applesa.ab.absxs.body_y\[5\] vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout761_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12701__B net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout859_A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_320_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09282__B game.CPU.applesa.ab.good_collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_4_clk_X clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16396__A net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_205_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10860_ _03499_ game.CPU.randy.counter1.count1\[14\] _03500_ game.CPU.randy.counter1.count1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__o22a_1
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09519_ net1102 net1269 vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_84_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_292_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09654__A1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10791_ _03342_ net561 vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__nor2_1
XANTENNA__09654__B2 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12429__A game.CPU.applesa.ab.absxs.body_x\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13024__S net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_234_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12530_ game.CPU.applesa.ab.absxs.body_x\[98\] net374 net527 game.CPU.applesa.ab.absxs.body_y\[97\]
+ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13738__A0 game.writer.tracker.frame\[209\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11052__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12461_ game.CPU.applesa.ab.absxs.body_y\[110\] net520 vssd1 vssd1 vccd1 vccd1 _06338_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_156_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_331_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_313_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13833__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14200_ game.CPU.applesa.ab.absxs.body_y\[67\] net945 vssd1 vssd1 vccd1 vccd1 _08074_
+ sky130_fd_sc_hd__xor2_1
X_11412_ game.CPU.applesa.ab.check_walls.above.walls\[115\] net762 vssd1 vssd1 vccd1
+ vccd1 _05301_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_340_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15180_ _03198_ _04580_ _03197_ vssd1 vssd1 vccd1 vccd1 _08756_ sky130_fd_sc_hd__a21oi_1
X_12392_ game.CPU.applesa.ab.absxs.body_x\[25\] net376 net369 _03350_ vssd1 vssd1
+ vccd1 vccd1 _06269_ sky130_fd_sc_hd__a22o_1
X_14131_ net1045 game.CPU.applesa.ab.check_walls.above.walls\[43\] vssd1 vssd1 vccd1
+ vccd1 _08005_ sky130_fd_sc_hd__xor2_1
X_11343_ net808 net259 net255 net809 _05231_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__o221a_1
XFILLER_0_132_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_278_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16152__B2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_238_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14163__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14062_ net1043 game.CPU.applesa.ab.check_walls.above.walls\[147\] vssd1 vssd1 vccd1
+ vccd1 _07936_ sky130_fd_sc_hd__xor2_1
XFILLER_0_293_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13505__A3 _07377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11274_ _04931_ _04932_ _04939_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_95_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_277_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13013_ game.writer.tracker.frame\[528\] game.writer.tracker.frame\[529\] net1007
+ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_245_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10225_ _04413_ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__or2_1
X_18870_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[0\] _00565_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__19732__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16455__A2 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17821_ _03148_ _03153_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__nor2_1
XANTENNA__09590__B1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18559__Q game.CPU.applesa.ab.absxs.body_y\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ net1260 _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_167_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold5 game.CPU.down_button.sync1.Q vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11508__A game.CPU.applesa.ab.check_walls.above.walls\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17752_ game.CPU.applesa.twoapples.count_luck\[0\] _03107_ _03109_ vssd1 vssd1 vccd1
+ vccd1 _03111_ sky130_fd_sc_hd__o21ai_1
X_10087_ _04293_ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__nor2_1
X_14964_ _08728_ _08733_ _08740_ vssd1 vssd1 vccd1 vccd1 _08741_ sky130_fd_sc_hd__or3b_1
X_16703_ _02484_ net63 _02567_ net1611 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[146\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_233_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11227__B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13915_ net984 game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1 vccd1
+ vccd1 _07789_ sky130_fd_sc_hd__xor2_1
XANTENNA__18936__D net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15922__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17683_ game.CPU.walls.rand_wall.count_luck\[3\] _03066_ vssd1 vssd1 vccd1 vccd1
+ _03068_ sky130_fd_sc_hd__and2_1
X_14895_ net1096 _08417_ vssd1 vssd1 vccd1 vccd1 _08672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19882__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload3_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19422_ clknet_leaf_43_clk game.writer.tracker.next_frame\[17\] net1306 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[17\] sky130_fd_sc_hd__dfrtp_1
X_16634_ net188 net124 _02391_ _02534_ net1468 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[110\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_334_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13846_ net281 _07713_ _07719_ net240 vssd1 vssd1 vccd1 vccd1 _07720_ sky130_fd_sc_hd__o211a_1
XFILLER_0_186_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19353_ clknet_leaf_71_clk _01363_ _00938_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.start_enable
+ sky130_fd_sc_hd__dfrtp_4
X_16565_ net1967 _02488_ _02490_ net127 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[85\]
+ sky130_fd_sc_hd__a22o_1
X_13777_ game.writer.tracker.frame\[149\] game.writer.tracker.frame\[151\] game.writer.tracker.frame\[152\]
+ game.writer.tracker.frame\[150\] net977 net1023 vssd1 vssd1 vccd1 vccd1 _07651_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__17168__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09645__A1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_256_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10989_ game.CPU.applesa.ab.absxs.body_x\[113\] net412 vssd1 vssd1 vccd1 vccd1 _04879_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__09645__B2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18304_ net641 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
X_15516_ _01499_ _01537_ _01492_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__a21boi_1
X_12728_ game.writer.tracker.frame\[98\] game.writer.tracker.frame\[99\] net995 vssd1
+ vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__mux2_1
X_19284_ clknet_leaf_68_clk _01333_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.enable
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16496_ net144 _02441_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__nor2_2
XANTENNA__16915__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_316_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12058__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18235_ net665 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
X_15447_ net879 _01473_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__or2_1
X_12659_ _03334_ game.CPU.applesa.twoapples.absxs.next_head\[6\] net361 game.CPU.applesa.ab.absxs.body_y\[64\]
+ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__a22o_1
XANTENNA__12626__X _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18026__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_303_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16472__C _02297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18166_ net610 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__inv_2
X_15378_ _08908_ _08912_ vssd1 vssd1 vccd1 vccd1 _08920_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12952__A1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19262__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17117_ _02365_ _02693_ net733 vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__o21a_1
Xhold405 game.CPU.kyle.L1.currentState\[5\] vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16143__A1 net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14329_ game.CPU.applesa.ab.absxs.body_x\[72\] net1072 vssd1 vssd1 vccd1 vccd1 _08203_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__09367__B game.CPU.applesa.ab.check_walls.above.walls\[34\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold416 game.writer.tracker.frame\[187\] vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
X_18097_ net634 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_345_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold427 game.writer.tracker.frame\[223\] vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold438 game.writer.tracker.frame\[461\] vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 game.writer.tracker.frame\[417\] vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
X_17048_ net188 _02412_ net91 _02685_ net1507 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[373\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__16694__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap179 net180 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_267_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ net1104 _03259_ game.CPU.applesa.ab.absxs.body_y\[108\] net893 _04112_ vssd1
+ vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__a221o_1
Xfanout907 _03199_ vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_209_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout918 _03194_ vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__buf_4
XANTENNA__10715__B1 _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout929 net930 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__buf_2
XANTENNA__16446__A2 _02243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18999_ net1194 _00226_ _00670_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[44\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12521__B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15654__B1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11137__B net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15832__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09884__A1 _03876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_356_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout175_A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10976__B net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_278_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout342_A game.CPU.walls.rand_wall.abduyd.next_wall\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09304_ net1132 game.CPU.applesa.ab.absxs.body_y\[55\] vssd1 vssd1 vccd1 vccd1 _03547_
+ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout1084_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12640__B1 game.CPU.applesa.twoapples.absxs.next_head\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_319_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13779__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09235_ game.CPU.applesa.ab.check_walls.above.walls\[193\] vssd1 vssd1 vccd1 vccd1
+ _03484_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19605__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_302_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout130_X net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10992__A game.CPU.applesa.ab.absxs.body_x\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13815__S0 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_X net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1251_A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1349_A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16921__A3 _02643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09166_ game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1 vccd1 vccd1
+ _03415_ sky130_fd_sc_hd__inv_2
XFILLER_0_302_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13291__S1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12943__A1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11746__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11600__B net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09097_ game.CPU.applesa.ab.absxs.body_y\[33\] vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1137_X net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_309_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09992__S _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19755__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13499__A2 _07073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout976_A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13367__X _07241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10706__B1 _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout88_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ net1163 game.CPU.applesa.out_random_2\[5\] vssd1 vssd1 vccd1 vccd1 _04218_
+ sky130_fd_sc_hd__nand2_2
XANTENNA__09293__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16437__A2 _02395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13527__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ game.CPU.apple_location\[0\] game.CPU.applesa.ab.apple_location\[0\] _04207_
+ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13019__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15742__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11047__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ game.CPU.applesa.ab.check_walls.above.walls\[68\] net394 _05847_ _05848_
+ _05201_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout931_X net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_240_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ game.writer.tracker.frame\[469\] game.writer.tracker.frame\[471\] game.writer.tracker.frame\[472\]
+ game.writer.tracker.frame\[470\] net975 net1014 vssd1 vssd1 vccd1 vccd1 _07574_
+ sky130_fd_sc_hd__mux4_1
X_10912_ _04807_ _04809_ _04257_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11615__X _05504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09740__B game.CPU.applesa.ab.check_walls.above.walls\[64\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19135__CLK net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10485__A2 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14680_ _08511_ _08512_ vssd1 vssd1 vccd1 vccd1 _08519_ sky130_fd_sc_hd__and2b_1
XANTENNA__13408__C1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11892_ net828 net303 _05775_ _05779_ _05354_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__o2111a_1
XANTENNA__14358__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13631_ game.writer.tracker.frame\[54\] net844 net838 game.writer.tracker.frame\[53\]
+ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10843_ _04743_ _04745_ _04742_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_211_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_343_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19003__Q game.CPU.applesa.ab.check_walls.above.walls\[48\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11063__A game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16350_ net134 net114 _02336_ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__or3_1
X_13562_ net220 _07423_ _07435_ net282 vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10774_ game.CPU.applesa.ab.absxs.body_y\[66\] _04679_ _04680_ game.CPU.applesa.ab.absxs.body_y\[62\]
+ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_181_Right_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19285__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15301_ game.CPU.applesa.twomode.number\[2\] _08844_ vssd1 vssd1 vccd1 vccd1 _08849_
+ sky130_fd_sc_hd__or2_1
X_12513_ _06383_ _06384_ _06388_ _06389_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__or4_1
X_16281_ net971 _02283_ _08028_ _06593_ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__14908__C1 game.CPU.applesa.ab.YMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_340_Left_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13493_ _07110_ _07112_ _07122_ _07111_ net700 net489 vssd1 vssd1 vccd1 vccd1 _07367_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18020_ net668 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12444_ game.CPU.applesa.ab.absxs.body_y\[106\] net520 net366 game.CPU.applesa.ab.absxs.body_y\[107\]
+ _06320_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__a221o_1
X_15232_ game.CPU.applesa.normal1.number\[2\] _08790_ game.CPU.applesa.normal1.counter
+ vssd1 vssd1 vccd1 vccd1 _08796_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_251_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12934__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11737__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15163_ net1214 net1239 net781 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__and3_1
XANTENNA__11510__B net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19450__RESET_B net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14524__D _08028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12375_ game.CPU.applesa.ab.absxs.body_x\[112\] net383 vssd1 vssd1 vccd1 vccd1 _06252_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14114_ _07986_ _07987_ vssd1 vssd1 vccd1 vccd1 _07988_ sky130_fd_sc_hd__nand2_1
X_11326_ net815 net316 vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__nor2_1
X_19971_ clknet_leaf_42_clk game.writer.tracker.next_frame\[566\] net1327 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[566\] sky130_fd_sc_hd__dfrtp_1
X_15094_ net1205 net1229 game.CPU.applesa.ab.check_walls.above.walls\[122\] vssd1
+ vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15917__B net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12147__C1 _06020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ net1053 game.CPU.applesa.ab.check_walls.above.walls\[194\] vssd1 vssd1 vccd1
+ vccd1 _07919_ sky130_fd_sc_hd__xor2_1
X_18922_ clknet_leaf_5_clk net1392 _00606_ vssd1 vssd1 vccd1 vccd1 game.CPU.left_button.eD1.Q1
+ sky130_fd_sc_hd__dfrtp_1
X_11257_ _05007_ _05008_ _05011_ _05016_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__or4_1
XANTENNA__14151__A3 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10208_ _04396_ _04397_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__nor2_1
X_18853_ clknet_leaf_6_clk _01244_ _00563_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.state\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_11188_ _03298_ net533 vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16979__A3 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_340_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17804_ net955 _03139_ _03140_ _01527_ vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__a22o_1
X_10139_ game.CPU.randy.f1.a1.count\[3\] game.CPU.randy.f1.a1.count\[2\] game.CPU.randy.f1.a1.count\[1\]
+ game.CPU.randy.f1.a1.count\[0\] vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__or4_1
X_18784_ clknet_leaf_11_clk _01201_ _00521_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[102\]
+ sky130_fd_sc_hd__dfrtp_4
X_15996_ _02003_ _02004_ _02005_ _02007_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09931__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15652__B net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17735_ game.CPU.applesa.ab.count\[0\] net1167 vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__nor2_1
X_14947_ game.CPU.walls.rand_wall.count_luck\[7\] game.CPU.walls.rand_wall.count_luck\[6\]
+ vssd1 vssd1 vccd1 vccd1 _08724_ sky130_fd_sc_hd__or2_1
XFILLER_0_221_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09650__B game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17666_ _03056_ net194 _03055_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__and3b_1
X_14878_ game.CPU.walls.abc.number\[2\] game.CPU.walls.abc.number\[6\] game.CPU.walls.abc.counter
+ vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19405_ clknet_leaf_47_clk game.writer.tracker.next_frame\[0\] net1294 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[0\] sky130_fd_sc_hd__dfrtp_1
X_16617_ net113 _02525_ net715 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__o21a_1
X_13829_ game.writer.tracker.frame\[542\] net842 net672 game.writer.tracker.frame\[544\]
+ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__o22a_1
XANTENNA__19628__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_253_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17597_ _03009_ _03014_ net585 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12069__A game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_327_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19336_ clknet_leaf_72_clk _01352_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.count_luck\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16548_ net1939 _02474_ _02478_ net129 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[80\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14555__Y game.CPU.walls.rand_wall.abduyd.next_wall\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_351_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19538__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13900__B net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19267_ clknet_leaf_8_clk _00055_ _00897_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_16479_ net169 _02348_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__and2_2
XFILLER_0_289_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16903__A3 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09020_ game.CPU.applesa.ab.absxs.body_x\[64\] vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__inv_2
XANTENNA__18652__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14375__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18218_ net666 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19778__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19198_ clknet_leaf_66_clk _01307_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.enable
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__16770__Y _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12516__B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11420__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18149_ net630 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__inv_2
Xhold202 game.writer.tracker.frame\[359\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_331_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold213 game.writer.tracker.frame\[480\] vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12616__C_N _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold224 game.writer.tracker.frame\[111\] vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14127__B1 game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold235 game.writer.tracker.frame\[381\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_348_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold246 game.writer.tracker.frame\[231\] vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15827__B net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14290__Y _08164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19008__CLK net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold257 game.writer.tracker.frame\[159\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15875__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold268 game.writer.tracker.frame\[526\] vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 game.writer.tracker.frame\[307\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _04148_ _04150_ _04151_ _04162_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__a31oi_1
XANTENNA__09825__B game.CPU.applesa.ab.absxs.body_x\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout704 net706 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout715 net717 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_113_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout726 _04738_ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_4
Xfanout737 net738 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_2
X_20042_ net1366 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_187_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09853_ _04094_ _04095_ _04092_ _04093_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__a211o_1
Xfanout748 net749 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12251__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout759 net760 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__buf_2
XANTENNA__17092__A2 _02486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_304_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15843__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ net1108 _03456_ game.CPU.applesa.ab.check_walls.above.walls\[146\] net920
+ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__a22o_1
XANTENNA__19158__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_283_Right_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_240_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10987__A game.CPU.applesa.ab.absxs.body_y\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13363__A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout557_A net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_202_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16674__A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout724_A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13650__X _07524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_X net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19961__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_315_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14194__A game.CPU.applesa.ab.absxs.body_x\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13169__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13302__S net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09218_ game.CPU.applesa.ab.check_walls.above.walls\[163\] vssd1 vssd1 vccd1 vccd1
+ _03467_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09288__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10490_ _04581_ _04612_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__nand2_1
XANTENNA__12426__B net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11719__A2 _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11330__B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09149_ game.CPU.applesa.ab.check_walls.above.walls\[35\] vssd1 vssd1 vccd1 vccd1
+ _03398_ sky130_fd_sc_hd__inv_2
XANTENNA__16107__B2 game.CPU.applesa.ab.absxs.body_y\[38\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14118__B1 game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16658__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12392__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12160_ game.CPU.applesa.ab.check_walls.above.walls\[39\] net296 net290 net822 vssd1
+ vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__a22o_1
XFILLER_0_258_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15737__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout881_X net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout979_X net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ game.CPU.applesa.ab.absxs.body_y\[34\] net541 vssd1 vssd1 vccd1 vccd1 _05001_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_92_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12091_ net804 net388 vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13341__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_290_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11042_ game.CPU.applesa.ab.absxs.body_y\[83\] net396 vssd1 vssd1 vccd1 vccd1 _04932_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_216_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17083__A2 _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15753__A _03381_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15850_ _03261_ net353 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_164_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16201__X _02213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14801_ game.CPU.randy.counter1.count\[8\] _08612_ net138 vssd1 vssd1 vccd1 vccd1
+ _08615_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_243_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_250_Right_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15781_ _01786_ _01792_ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__or2_1
XANTENNA__09848__A1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13644__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ game.writer.tracker.frame\[562\] game.writer.tracker.frame\[563\] net1021
+ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09848__B2 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17520_ game.CPU.modea.Qa\[0\] _02849_ _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__a21o_1
XFILLER_0_231_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11655__A1 game.CPU.applesa.ab.check_walls.above.walls\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14732_ _08561_ _08562_ net54 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__and3b_1
X_11944_ net796 net310 vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__or2_1
X_17451_ net1459 net264 _02869_ _02880_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_318_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11875_ game.CPU.applesa.ab.check_walls.above.walls\[143\] net310 vssd1 vssd1 vccd1
+ vccd1 _05763_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14663_ _08491_ _08501_ vssd1 vssd1 vccd1 vccd1 _08502_ sky130_fd_sc_hd__and2_1
XFILLER_0_345_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16402_ net115 net164 net68 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13614_ _07475_ _07479_ _07483_ _07487_ net244 vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_45_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ _04482_ _04568_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__or2_1
XANTENNA__18675__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_253_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12604__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17382_ _02792_ _02802_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__nand2_1
X_14594_ game.CPU.clock1.counter\[1\] game.CPU.clock1.counter\[0\] game.CPU.clock1.counter\[2\]
+ vssd1 vssd1 vccd1 vccd1 _08454_ sky130_fd_sc_hd__a21o_1
XANTENNA__19920__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19121_ net1182 _00161_ _00792_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[166\]
+ sky130_fd_sc_hd__dfrtp_1
X_16333_ game.writer.tracker.frame\[20\] net735 _02323_ vssd1 vssd1 vccd1 vccd1 _02324_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13545_ _07412_ _07416_ net226 vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10757_ game.CPU.applesa.ab.absxs.body_y\[99\] net263 _04719_ game.CPU.applesa.ab.absxs.body_y\[95\]
+ vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_175_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19052_ net1191 _00284_ _00723_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[97\]
+ sky130_fd_sc_hd__dfrtp_4
X_13476_ _07152_ _07154_ net700 vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__mux2_1
X_16264_ _02230_ _02268_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__or2_2
XANTENNA__16897__A2 _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_353_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ game.CPU.applesa.ab.absxs.body_y\[101\] _04595_ _04708_ game.CPU.applesa.ab.absxs.body_y\[97\]
+ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18003_ net634 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__inv_2
XANTENNA__11240__B net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15215_ net758 _08778_ _08779_ _08780_ _08781_ vssd1 vssd1 vccd1 vccd1 _08782_ sky130_fd_sc_hd__a32o_1
X_12427_ game.CPU.applesa.ab.absxs.body_y\[103\] net367 vssd1 vssd1 vccd1 vccd1 _06304_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_298_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15928__A _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16195_ _01626_ _01630_ _01631_ _01633_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__or4_1
XFILLER_0_341_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16649__A2 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13580__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ game.CPU.applesa.ab.absxs.body_x\[44\] net383 vssd1 vssd1 vccd1 vccd1 _06235_
+ sky130_fd_sc_hd__xnor2_1
X_15146_ net1213 net1240 game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1
+ vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__and3_1
XANTENNA__10394__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10394__B2 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11309_ game.CPU.applesa.ab.check_walls.above.walls\[67\] net763 vssd1 vssd1 vccd1
+ vccd1 _05198_ sky130_fd_sc_hd__xor2_2
X_19954_ clknet_leaf_43_clk game.writer.tracker.next_frame\[549\] net1303 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[549\] sky130_fd_sc_hd__dfrtp_1
X_15077_ net1212 net1238 game.CPU.applesa.ab.check_walls.above.walls\[105\] vssd1
+ vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__and3_1
X_12289_ net830 net549 vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__and2_1
XANTENNA__12352__A game.CPU.applesa.ab.absxs.body_y\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_266_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_264_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13332__A1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14028_ net1069 _03464_ _03467_ net1043 vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__a22o_1
XANTENNA__09536__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18905_ clknet_leaf_4_clk _01272_ _00589_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_19885_ clknet_leaf_27_clk game.writer.tracker.next_frame\[480\] net1311 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[480\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_206_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11343__B1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17074__A2 _02693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18836_ clknet_leaf_0_clk _01227_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10697__A2 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18767_ clknet_leaf_50_clk _01184_ _00504_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[69\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09839__A1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15979_ game.CPU.applesa.ab.check_walls.above.walls\[66\] net468 vssd1 vssd1 vccd1
+ vccd1 _01991_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_334_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13635__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19450__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09839__B2 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17718_ game.CPU.applesa.ab.count_luck\[2\] game.CPU.applesa.ab.count_luck\[1\] _03086_
+ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__and3_1
X_18698_ clknet_leaf_12_clk _01115_ _00435_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[48\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_353_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_348_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17649_ game.CPU.kyle.L1.cnt_500hz\[7\] _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__or2_1
XANTENNA__11415__B net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_44_clk_X clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16585__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16494__A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_275_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13494__S1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17129__A3 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19319_ clknet_leaf_71_clk _01343_ _00925_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.apple_location2_n\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16337__A1 net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_317_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12527__A game.CPU.applesa.ab.absxs.body_y\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11431__A game.CPU.applesa.ab.check_walls.above.walls\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_59_clk_X clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13246__S1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09003_ game.CPU.applesa.ab.absxs.body_x\[107\] vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__inv_2
XANTENNA__12246__B net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10047__A net1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout305_A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1047_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09395__X _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__B1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_257_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_352_Right_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_306_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15848__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12262__A net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13859__C1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_228_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1214_A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout512 net514 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12757__S0 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ game.CPU.bodymain1.Direction\[0\] net1261 vssd1 vssd1 vccd1 vccd1 _04147_
+ sky130_fd_sc_hd__and2b_1
Xfanout523 net527 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_4
Xfanout534 net537 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_4
XANTENNA_fanout674_A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_X net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 net546 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_4
Xfanout556 net557 vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_4
XANTENNA__17065__A2 _02449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_272_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20025_ net1276 vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_09836_ net927 game.CPU.applesa.ab.absxs.body_x\[107\] _03254_ net1102 _04076_ vssd1
+ vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__o221a_1
XANTENNA__09842__Y _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout567 net568 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_4
Xfanout578 net579 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_4
Xfanout589 net590 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_2
XANTENNA__16388__B net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16273__B1 _02267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16812__A2 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ net1155 _03433_ game.CPU.applesa.ab.check_walls.above.walls\[102\] net903
+ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_244_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14189__A game.CPU.applesa.ab.absxs.body_y\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12834__A0 _06704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18698__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09698_ _03931_ _03935_ _03938_ _03940_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__or4_2
XFILLER_0_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19943__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_317_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11325__B net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13821__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11660_ _03385_ _05194_ _05206_ _05547_ _05548_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__o311a_1
XFILLER_0_193_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_354_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10611_ game.CPU.applesa.ab.absxs.body_x\[80\] _04673_ _04674_ net1267 vssd1 vssd1
+ vccd1 vccd1 _01131_ sky130_fd_sc_hd__a22o_1
X_11591_ game.CPU.applesa.ab.check_walls.above.walls\[105\] net770 vssd1 vssd1 vccd1
+ vccd1 _05480_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_354_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12437__A game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_289_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13330_ _06704_ _06741_ _06742_ _06743_ net500 net695 vssd1 vssd1 vccd1 vccd1 _07204_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_107_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10542_ game.CPU.applesa.ab.absxs.body_x\[38\] _04642_ _04643_ game.CPU.applesa.ab.absxs.body_x\[34\]
+ vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_340_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12156__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13261_ game.writer.tracker.frame\[488\] game.writer.tracker.frame\[489\] net1000
+ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__mux2_1
XANTENNA__15748__A game.CPU.applesa.ab.check_walls.above.walls\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11060__B net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10473_ net929 game.CPU.applesa.ab.absxs.body_x\[90\] vssd1 vssd1 vccd1 vccd1 _04603_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_323_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12365__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19323__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12212_ game.CPU.applesa.ab.check_walls.above.walls\[174\] net418 vssd1 vssd1 vccd1
+ vccd1 _06098_ sky130_fd_sc_hd__xnor2_1
X_15000_ net1223 net1251 net826 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__and3_1
XFILLER_0_350_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13562__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_328_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13192_ game.writer.tracker.frame\[408\] game.writer.tracker.frame\[409\] net1036
+ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10376__A1 net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10376__B2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ game.CPU.applesa.ab.check_walls.above.walls\[189\] net386 vssd1 vssd1 vccd1
+ vccd1 _06030_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_349_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_248_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16951_ _02398_ net93 _02656_ game.writer.tracker.frame\[305\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[305\] sky130_fd_sc_hd__a22o_1
X_12074_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__inv_2
XFILLER_0_263_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19473__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_285_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17056__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13555__X _07429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ game.CPU.applesa.ab.absxs.body_y\[90\] net403 vssd1 vssd1 vccd1 vccd1 _04915_
+ sky130_fd_sc_hd__nand2_1
X_15902_ _01904_ _01905_ _01911_ _01912_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a22o_1
X_19670_ clknet_leaf_32_clk game.writer.tracker.next_frame\[265\] net1292 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[265\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_218_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10679__A2 game.CPU.applesa.ab.absxs.body_x\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_263_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16882_ net177 net135 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__nand2_4
XANTENNA__11876__B2 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18621_ clknet_leaf_13_clk _01038_ _00358_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[115\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16803__A2 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15833_ game.CPU.applesa.ab.absxs.body_x\[108\] net272 vssd1 vssd1 vccd1 vccd1 _01845_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_189_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18567__Q game.CPU.applesa.ab.absxs.body_y\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_263_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09912__C net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18552_ clknet_leaf_45_clk _00975_ net1298 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.cmd_num\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11628__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15764_ game.CPU.applesa.ab.absxs.body_x\[118\] net467 vssd1 vssd1 vccd1 vccd1 _01776_
+ sky130_fd_sc_hd__xnor2_1
X_12976_ net488 _06849_ _06848_ net228 vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__o211a_1
X_17503_ game.CPU.luck1.Qa\[0\] _02774_ net428 _02860_ vssd1 vssd1 vccd1 vccd1 _02932_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11235__B net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14715_ _03511_ _08549_ vssd1 vssd1 vccd1 vccd1 _08551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_358_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_346_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19812__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15930__B net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11927_ net748 _05507_ _05511_ _05512_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__o211a_1
X_18483_ net638 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__inv_2
X_15695_ _03315_ net336 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13290__X _07164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_345_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17434_ net1124 _02784_ _02824_ _02830_ _02863_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__a2111o_1
X_14646_ net741 _08451_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_body_clk sky130_fd_sc_hd__and2_1
XFILLER_0_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_318_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11858_ net751 _05490_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_345_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_19 _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17365_ _03196_ _02789_ _02791_ _02794_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__o31ai_1
XANTENNA__12053__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ game.CPU.applesa.ab.absxs.body_y\[16\] _04699_ _04700_ game.CPU.applesa.ab.absxs.body_y\[12\]
+ vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__a22o_1
XFILLER_0_172_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14577_ game.CPU.clock1.counter\[17\] game.CPU.clock1.counter\[20\] vssd1 vssd1 vccd1
+ vccd1 _08439_ sky130_fd_sc_hd__nand2_1
XANTENNA__12053__B2 game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ net570 _05253_ net395 game.CPU.applesa.ab.check_walls.above.walls\[36\] _05676_
+ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19104_ net1180 _00142_ _00775_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[149\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_172_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16316_ _02273_ _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ game.writer.tracker.frame\[93\] game.writer.tracker.frame\[95\] game.writer.tracker.frame\[96\]
+ game.writer.tracker.frame\[94\] net976 net1017 vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__mux4_1
XANTENNA__10603__A2 _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17296_ net2050 net721 _02755_ _02374_ net175 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[551\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_250_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12066__B net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__A1_N net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19035_ net1191 _00266_ _00706_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[80\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12781__S net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16247_ _02228_ _02253_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__or2_1
XANTENNA__15658__A game.CPU.applesa.ab.check_walls.above.walls\[48\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13459_ net496 _07332_ _07331_ net230 vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__a211o_1
XANTENNA__15542__A2 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18034__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16106__X _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_212_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_301_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_71_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16178_ _02026_ _02028_ _02131_ _02189_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__or4_4
XANTENNA__10367__A1 game.CPU.applesa.ab.absxs.body_y\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14281__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19816__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09375__B game.CPU.applesa.ab.check_walls.above.walls\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15129_ net1208 net1234 game.CPU.applesa.ab.check_walls.above.walls\[157\] vssd1
+ vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15096__C game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_282_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19937_ clknet_leaf_42_clk game.writer.tracker.next_frame\[532\] net1326 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[532\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16489__A net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_184_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17047__A2 _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13906__A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19868_ clknet_leaf_20_clk game.writer.tracker.next_frame\[463\] net1308 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[463\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11867__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_345_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19966__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11405__A1_N net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13069__A0 game.writer.tracker.frame\[200\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_301_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09621_ net1112 game.CPU.applesa.ab.check_walls.above.walls\[0\] vssd1 vssd1 vccd1
+ vccd1 _03864_ sky130_fd_sc_hd__xor2_1
X_18819_ clknet_leaf_73_clk game.CPU.clock1.next_body_clk _00556_ vssd1 vssd1 vccd1
+ vccd1 game.CPU.applesa.clk_body sky130_fd_sc_hd__dfrtp_2
X_19799_ clknet_leaf_33_clk game.writer.tracker.next_frame\[394\] net1328 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[394\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13117__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ net1087 game.CPU.applesa.ab.absxs.body_x\[115\] vssd1 vssd1 vccd1 vccd1 _03795_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__11426__A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_223_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10330__A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09483_ net915 game.CPU.applesa.ab.check_walls.above.walls\[177\] game.CPU.applesa.ab.check_walls.above.walls\[178\]
+ net921 _03725_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__o221a_1
XANTENNA__11145__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15840__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12956__S net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout255_A _05207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18209__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14456__B net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_195_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_24_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_336_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout422_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12257__A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_351_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19346__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_312_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12595__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10048__Y _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_X net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14472__A game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_171_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_305_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13544__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12347__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_277_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14191__B net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19496__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_A _03368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17286__A2 _02258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_319_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1307 net1360 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__buf_2
Xfanout320 game.CPU.applesa.ab.absxs.next_head\[2\] vssd1 vssd1 vccd1 vccd1 net320
+ sky130_fd_sc_hd__buf_4
Xfanout1318 net1323 vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__buf_2
XFILLER_0_245_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1329 net1333 vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__clkbuf_4
Xfanout342 game.CPU.walls.rand_wall.abduyd.next_wall\[4\] vssd1 vssd1 vccd1 vccd1
+ net342 sky130_fd_sc_hd__buf_6
Xfanout353 game.CPU.walls.rand_wall.abduyd.next_wall\[1\] vssd1 vssd1 vccd1 vccd1
+ net353 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_148_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_323_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12720__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout364 net368 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_255_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout375 _06209_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_8
X_20008_ net1377 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_161_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09819_ net924 game.CPU.applesa.ab.absxs.body_x\[27\] _03279_ net1091 vssd1 vssd1
+ vccd1 vccd1 _04062_ sky130_fd_sc_hd__a22o_1
Xfanout397 net400 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_4
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11251__A2_N net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10530__B2 game.CPU.applesa.ab.absxs.body_x\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11336__A game.CPU.applesa.ab.check_walls.above.walls\[80\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12830_ game.writer.tracker.frame\[288\] game.writer.tracker.frame\[289\] net1001
+ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__mux2_2
XFILLER_0_201_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15750__B net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_328_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16549__A1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12761_ _06581_ _06586_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__and2_1
XFILLER_0_213_298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_295_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16549__B2 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14500_ game.CPU.apple_location\[5\] net958 vssd1 vssd1 vccd1 vccd1 _08374_ sky130_fd_sc_hd__or2_1
XFILLER_0_327_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17210__A2 net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ game.CPU.applesa.ab.apple_possible\[7\] _05599_ vssd1 vssd1 vccd1 vccd1 _05600_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_237_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _06554_ _06565_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__nand2_1
X_15480_ _08925_ _08931_ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__or2_2
XFILLER_0_68_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ game.CPU.applesa.ab.check_walls.above.walls\[156\] net249 vssd1 vssd1 vccd1
+ vccd1 _05532_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14431_ game.CPU.applesa.ab.absxs.body_x\[24\] net887 net1045 _03278_ vssd1 vssd1
+ vccd1 vccd1 _08305_ sky130_fd_sc_hd__a22o_1
XFILLER_0_343_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_351_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16862__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12167__A game.CPU.applesa.ab.check_walls.above.walls\[157\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_315_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17150_ _02425_ _02693_ net737 vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__o21a_1
XFILLER_0_181_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ net742 _05460_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14362_ game.CPU.applesa.ab.absxs.body_x\[100\] net1072 vssd1 vssd1 vccd1 vccd1 _08236_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_172_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11794__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16101_ _03353_ net339 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__xnor2_1
X_13313_ net224 _07186_ _07185_ net274 vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__a211o_1
X_10525_ _04636_ game.CPU.applesa.ab.absxs.body_x\[60\] _04632_ vssd1 vssd1 vccd1
+ vccd1 _01179_ sky130_fd_sc_hd__mux2_1
XANTENNA__19839__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17081_ _02300_ net57 _02696_ net1808 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[395\]
+ sky130_fd_sc_hd__a22o_1
X_14293_ game.CPU.applesa.ab.absxs.body_y\[55\] net946 vssd1 vssd1 vccd1 vccd1 _08167_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_220_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13244_ game.writer.tracker.frame\[502\] game.writer.tracker.frame\[503\] net1015
+ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__mux2_1
X_16032_ _02040_ _02041_ _02042_ _02043_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__or4_1
XANTENNA__09476__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10456_ _04358_ _04579_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__nor2_4
XFILLER_0_220_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ game.writer.tracker.frame\[444\] game.writer.tracker.frame\[445\] net1038
+ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_248_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10387_ net1153 game.CPU.apple_location\[4\] vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_290_Left_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16485__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19989__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18863__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ _05397_ _05399_ _05400_ _05402_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__or4b_1
XANTENNA__13299__A0 _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_264_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_261_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17983_ net606 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__inv_2
X_19722_ clknet_leaf_35_clk game.writer.tracker.next_frame\[317\] net1346 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[317\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17029__A2 _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16934_ net184 _02524_ net87 _02651_ net1599 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[293\]
+ sky130_fd_sc_hd__a32o_1
X_12057_ _05442_ _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__nand2_1
XANTENNA__16102__A game.CPU.applesa.ab.absxs.body_y\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11008_ _03306_ net401 vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__nor2_1
XANTENNA_output51_A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19653_ clknet_leaf_22_clk game.writer.tracker.next_frame\[248\] net1343 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[248\] sky130_fd_sc_hd__dfrtp_1
X_16865_ net133 _02418_ net123 _02626_ net1876 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[248\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__16788__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18604_ clknet_leaf_3_clk _00006_ _00341_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.row_2\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_15816_ _03264_ net269 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__xnor2_1
X_19584_ clknet_leaf_35_clk game.writer.tracker.next_frame\[179\] net1338 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[179\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16252__A3 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16796_ _02473_ net98 net716 vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__o21a_1
XANTENNA__14263__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18535_ net611 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__inv_2
XFILLER_0_204_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15747_ _03380_ net334 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15660__B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ net217 _06778_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__and2_1
XANTENNA__13471__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_259_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19369__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18466_ net652 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__inv_2
X_15678_ _03382_ net271 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_272_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17417_ _03217_ game.CPU.kyle.L1.nextState\[2\] _02816_ vssd1 vssd1 vccd1 vccd1 _02847_
+ sky130_fd_sc_hd__or3_2
X_14629_ game.CPU.clock1.counter\[15\] _08474_ net267 vssd1 vssd1 vccd1 vccd1 _08476_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_346_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_261_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18397_ net617 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__inv_2
XANTENNA__16960__A1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_333_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17348_ net1258 _03219_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__nor2_4
XFILLER_0_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12982__C1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18760__Q game.CPU.applesa.ab.absxs.body_x\[54\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17279_ net117 _02574_ _02750_ net1956 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[539\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_348_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12329__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09386__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19018_ net1196 _00247_ _00689_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12524__B net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_302_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17268__A2 _02322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15835__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ game.CPU.applesa.ab.absxs.body_x\[86\] vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__inv_2
XANTENNA__13829__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_225_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10760__A1 game.CPU.applesa.ab.absxs.body_y\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_299_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_282_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10612__X _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10979__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout372_A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15851__A game.CPU.applesa.ab.absxs.body_x\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09604_ _03841_ _03842_ _03843_ _03846_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__or4_1
XFILLER_0_155_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16666__B _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_197_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11068__A2 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09535_ net911 game.CPU.applesa.ab.check_walls.above.walls\[72\] _03422_ net1156
+ _03777_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout160_X net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10995__A game.CPU.applesa.ab.absxs.body_y\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1281_A net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11989__A1_N game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_X net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09466_ game.CPU.applesa.ab.absxs.body_y\[92\] net892 net1136 _03296_ vssd1 vssd1
+ vccd1 vccd1 _03709_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10815__A2 game.CPU.applesa.ab.absxs.body_y\[113\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18736__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11603__B net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09397_ net1110 game.CPU.applesa.ab.check_walls.above.walls\[88\] vssd1 vssd1 vccd1
+ vccd1 _03640_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16951__A1 _02398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16951__B2 game.writer.tracker.frame\[305\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09995__S _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18670__Q game.CPU.applesa.ab.absxs.body_y\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16703__A1 _02484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1334_X net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13517__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10310_ game.CPU.randy.f1.a1.count\[9\] _04491_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__and2_1
XANTENNA__18886__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11290_ _05140_ _05179_ _05178_ _04962_ _05084_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_131_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__Y _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_325_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17259__A2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ _04415_ _04431_ _04432_ _04433_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15585__X _01597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18402__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_18_Left_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12740__A2 _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ net1134 _04362_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout961_X net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15745__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10751__A1 game.CPU.applesa.ab.absxs.body_y\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1104 game.CPU.applesa.ab.snake_head_x\[1\] vssd1 vssd1 vccd1 vccd1 net1104
+ sky130_fd_sc_hd__buf_4
Xfanout1115 game.CPU.bodymain1.main.score\[5\] vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__buf_2
Xfanout1126 net1129 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09743__B game.CPU.applesa.ab.check_walls.above.walls\[70\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14980_ net1225 net1252 game.CPU.applesa.ab.check_walls.above.walls\[8\] vssd1 vssd1
+ vccd1 vccd1 _00165_ sky130_fd_sc_hd__and3_1
Xfanout1137 net1138 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12450__A game.CPU.applesa.ab.absxs.body_x\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout150 net151 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_218_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1148 net1151 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__clkbuf_8
Xfanout161 _02256_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_273_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1159 net1160 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__buf_4
Xfanout172 _02254_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_89_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout183 net184 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_4
X_13931_ net961 net823 vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__nand2_1
Xfanout194 _03037_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09462__C net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19006__Q game.CPU.applesa.ab.check_walls.above.walls\[51\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10503__A1 game.CPU.applesa.ab.absxs.body_x\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_282_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10503__B2 game.CPU.applesa.ab.absxs.body_x\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16650_ net190 net128 _02412_ _02543_ net1760 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[117\]
+ sky130_fd_sc_hd__a32o_1
X_13862_ game.writer.tracker.frame\[550\] net842 net835 game.writer.tracker.frame\[549\]
+ net274 vssd1 vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__o221a_1
XFILLER_0_159_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19511__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16576__B _02376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15601_ game.CPU.applesa.ab.check_walls.above.walls\[112\] net354 vssd1 vssd1 vccd1
+ vccd1 _01613_ sky130_fd_sc_hd__xnor2_1
X_12813_ _06683_ _06686_ net678 vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16581_ net1692 _02500_ _02501_ net126 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[90\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_241_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13793_ net215 _07666_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_27_Left_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18320_ net615 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__inv_2
X_15532_ _06562_ _01551_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12744_ _06569_ _06577_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10806__A2 _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14096__B net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18251_ net622 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_328_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15463_ _01432_ _01440_ _01481_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__nor3_1
XFILLER_0_60_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11513__B net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19661__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16942__A1 _02299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ net1075 net1057 vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__nor2_1
XFILLER_0_343_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17202_ _02513_ net71 _02731_ net1872 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[481\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_181_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12559__A2 game.CPU.applesa.twoapples.absxs.next_head\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14414_ game.CPU.applesa.ab.absxs.body_x\[45\] net884 net878 game.CPU.applesa.ab.absxs.body_x\[46\]
+ vssd1 vssd1 vccd1 vccd1 _08288_ sky130_fd_sc_hd__a22o_1
X_11626_ net742 _05507_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__xnor2_1
X_18182_ net610 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__inv_2
X_15394_ _03363_ game.writer.updater.commands.mode\[0\] vssd1 vssd1 vccd1 vccd1 _08936_
+ sky130_fd_sc_hd__nand2_2
XANTENNA__09424__A2 game.CPU.applesa.ab.check_walls.above.walls\[115\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17133_ net165 net67 net76 _02712_ net1532 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[431\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14345_ _03246_ net1072 net987 _03313_ _08215_ vssd1 vssd1 vccd1 vccd1 _08219_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11557_ net743 _05441_ _05443_ _05444_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__o211a_1
XANTENNA__13508__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_330_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17064_ _02438_ _02455_ _02689_ net1913 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[385\]
+ sky130_fd_sc_hd__a22o_1
Xhold609 game.writer.tracker.frame\[537\] vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
X_10508_ game.CPU.applesa.ab.absxs.body_x\[71\] _04625_ _04626_ game.CPU.applesa.ab.absxs.body_x\[67\]
+ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__a22o_1
X_14276_ game.CPU.applesa.ab.absxs.body_x\[50\] net880 net985 _03342_ _08149_ vssd1
+ vssd1 vccd1 vccd1 _08150_ sky130_fd_sc_hd__o221a_1
X_11488_ _05362_ _05363_ _05376_ _05361_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__a31o_1
XANTENNA__16170__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12344__B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16015_ _03477_ net343 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10497__D_N net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14181__A1 game.CPU.applesa.ab.absxs.body_x\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13227_ _07099_ _07100_ net498 vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__mux2_1
X_10439_ net1966 net847 _04165_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__a21o_1
XANTENNA__14181__B2 game.CPU.applesa.ab.absxs.body_y\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_249_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18312__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ game.writer.tracker.frame\[160\] game.writer.tracker.frame\[161\] net1023
+ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__mux2_2
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15655__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19041__CLK net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ _05364_ _05365_ _05369_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__nand3_1
X_13089_ net700 _06962_ _06959_ net209 vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__o211a_1
XFILLER_0_264_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17966_ net668 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__inv_2
XANTENNA__12360__A game.CPU.applesa.ab.absxs.body_x\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09653__B game.CPU.applesa.ab.check_walls.above.walls\[171\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18609__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_181_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16917_ _02497_ net95 _02647_ net1818 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[280\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_251_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19705_ clknet_leaf_31_clk game.writer.tracker.next_frame\[300\] net1284 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[300\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13692__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17897_ net643 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__inv_2
XFILLER_0_192_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16848_ net1464 _02620_ _02621_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[237\]
+ sky130_fd_sc_hd__a21o_1
X_19636_ clknet_leaf_28_clk game.writer.tracker.next_frame\[231\] net1287 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[231\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19191__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_195_Right_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_220_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14558__Y game.CPU.walls.rand_wall.abduyd.next_wall\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18755__Q game.CPU.applesa.ab.absxs.body_x\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19567_ clknet_leaf_48_clk game.writer.tracker.next_frame\[162\] net1296 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[162\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18759__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13903__B net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16779_ _02445_ net99 net730 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__o21a_1
XFILLER_0_342_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13191__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09320_ net1103 game.CPU.applesa.ab.absxs.body_x\[65\] vssd1 vssd1 vccd1 vccd1 _03563_
+ sky130_fd_sc_hd__xor2_1
X_18518_ net588 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17186__A1 _02490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19498_ clknet_leaf_25_clk game.writer.tracker.next_frame\[93\] net1321 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[93\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12519__B net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_307_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09251_ game.CPU.randy.counter1.count\[14\] vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__inv_2
X_18449_ net592 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__inv_2
XANTENNA__11470__A2 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16933__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_192_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09182_ game.CPU.applesa.ab.check_walls.above.walls\[96\] vssd1 vssd1 vccd1 vccd1
+ _03431_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11758__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14023__A2_N net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout120_A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09828__B game.CPU.applesa.ab.absxs.body_x\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13130__S net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_314_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_299_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_231_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12254__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1127_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17110__A1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10733__A1 game.CPU.applesa.ab.absxs.body_y\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10733__B2 game.CPU.applesa.ab.absxs.body_y\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16464__A3 _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ game.CPU.applesa.ab.absxs.body_y\[7\] vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__inv_2
XANTENNA__19534__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14475__A2 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_320_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13683__A0 game.writer.tracker.frame\[449\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout754_A _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_316_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_316_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout921_A _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19684__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19203__D _00016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_357_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09518_ net1102 net1269 vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10790_ net937 game.CPU.applesa.ab.absxs.body_y\[45\] net562 _04726_ vssd1 vssd1
+ vccd1 vccd1 _01004_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_292_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12429__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11997__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_234_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09449_ net925 game.CPU.applesa.ab.check_walls.above.walls\[139\] _03454_ net1145
+ _03687_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__o221a_1
XANTENNA__16924__A1 _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14484__X _08358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17301__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12460_ game.CPU.applesa.ab.absxs.body_x\[108\] net382 vssd1 vssd1 vccd1 vccd1 _06337_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_331_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11749__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_313_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11411_ net796 net259 vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__nor2_1
XANTENNA__12410__A1 game.CPU.applesa.ab.absxs.body_x\[53\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12391_ game.CPU.applesa.ab.absxs.body_x\[26\] net374 vssd1 vssd1 vccd1 vccd1 _06268_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_352_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11342_ _04460_ _05223_ _05226_ net743 _05230_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__o221a_1
X_14130_ net1054 game.CPU.applesa.ab.check_walls.above.walls\[42\] vssd1 vssd1 vccd1
+ vccd1 _08004_ sky130_fd_sc_hd__xor2_1
XFILLER_0_278_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_278_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16152__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19064__CLK net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14163__A1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14163__B2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11273_ _04933_ _04934_ _04935_ _04937_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__or4_1
X_14061_ _07928_ _07929_ _07933_ _07934_ vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__a211o_1
XANTENNA__15756__A game.CPU.applesa.ab.absxs.body_x\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_238_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_297_Right_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13012_ game.writer.tracker.frame\[520\] game.writer.tracker.frame\[521\] net1005
+ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__mux2_1
XANTENNA__09754__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _04373_ _04388_ _04412_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_37_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19656__RESET_B net1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_245_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10724__A1 game.CPU.applesa.ab.absxs.body_y\[38\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10724__B2 game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13349__S0 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17820_ game.writer.updater.commands.count\[2\] game.writer.updater.commands.count\[1\]
+ game.writer.updater.commands.count\[0\] vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__and3_1
XANTENNA__09590__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17971__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ game.CPU.randy.f1.state\[1\] game.CPU.randy.f1.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _04350_ sky130_fd_sc_hd__nand2_1
XANTENNA__09590__B2 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16455__A3 _02412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14466__A2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15663__B2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17751_ game.CPU.applesa.twoapples.count_luck\[0\] _03107_ vssd1 vssd1 vccd1 vccd1
+ _03110_ sky130_fd_sc_hd__and2_1
XFILLER_0_261_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6 game.CPU.reset_button1.sync1.Q vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ _04288_ _04292_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__xnor2_1
X_14963_ _08665_ _08735_ _08738_ _08739_ vssd1 vssd1 vccd1 vccd1 _08740_ sky130_fd_sc_hd__o211a_1
XANTENNA__11508__B net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16702_ _02482_ net63 _02567_ net1660 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[145\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15491__A _08027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18901__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13914_ _07784_ _07785_ _07786_ _07787_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__or4_1
XANTENNA__09342__B2 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17682_ _03062_ _03066_ _03067_ vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__nor3_1
X_14894_ net1096 _08417_ vssd1 vssd1 vccd1 vccd1 _08671_ sky130_fd_sc_hd__nand2_1
X_19421_ clknet_leaf_43_clk game.writer.tracker.next_frame\[16\] net1303 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[16\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16612__B1 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16633_ _02389_ _02518_ _02534_ net1613 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[109\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_226_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13845_ net506 _07716_ _07717_ _07718_ net275 vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__a311o_1
XFILLER_0_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19352_ net1167 _01362_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.normal1.counter_flip
+ sky130_fd_sc_hd__dfxtp_1
X_16564_ net154 _02489_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__and2_1
X_13776_ net512 _07645_ _07646_ _07649_ vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__a31o_1
XANTENNA__17168__A1 _02462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_256_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10988_ _03323_ game.CPU.applesa.ab.absxs.next_head\[5\] vssd1 vssd1 vccd1 vccd1
+ _04878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11988__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18303_ net643 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
X_15515_ _01434_ _01490_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__nand2_1
XANTENNA__11243__B net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12727_ game.writer.tracker.frame\[104\] game.writer.tracker.frame\[105\] net995
+ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__mux2_1
X_19283_ clknet_leaf_68_clk _01332_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.count\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_356_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_316_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16495_ _08404_ _01515_ _02357_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_178_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_328_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18234_ net665 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__inv_2
X_15446_ net1076 net1065 net1048 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__o21ai_1
X_12658_ _06373_ _06534_ _06374_ _06533_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__or4b_1
XFILLER_0_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12456__A2_N net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19407__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11609_ game.CPU.applesa.ab.check_walls.above.walls\[100\] net253 net316 net804 vssd1
+ vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__a2bb2o_1
X_18165_ net629 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__inv_2
X_15377_ _08918_ vssd1 vssd1 vccd1 vccd1 _08919_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12589_ net1268 net528 net359 game.CPU.applesa.ab.absxs.body_y\[88\] _06465_ vssd1
+ vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__o221a_1
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Left_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_10_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
X_17116_ _02364_ net80 _02706_ net1982 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[419\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14328_ game.CPU.applesa.ab.absxs.body_x\[72\] net1072 vssd1 vssd1 vccd1 vccd1 _08202_
+ sky130_fd_sc_hd__or2_1
X_18096_ net605 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__inv_2
Xhold406 game.writer.tracker.frame\[444\] vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16143__A2 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_345_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_296_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold417 game.writer.tracker.frame\[535\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_187_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold428 game.writer.tracker.frame\[523\] vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17047_ net188 _02410_ net91 _02685_ net1503 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[372\]
+ sky130_fd_sc_hd__a32o_1
Xhold439 game.writer.tracker.frame\[517\] vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14259_ game.CPU.applesa.ab.absxs.body_y\[79\] net941 vssd1 vssd1 vccd1 vccd1 _08133_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19557__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_267_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_264_Right_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09664__A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13901__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 net909 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_209_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10715__B2 game.CPU.applesa.ab.absxs.body_y\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout919 net921 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11912__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09581__A1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16446__A3 _02405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__B2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18998_ net1195 _00225_ _00669_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[43\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_209_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17949_ net613 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__inv_2
XANTENNA__18581__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_240_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Left_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16603__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09884__A2 _03880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_356_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19619_ clknet_leaf_21_clk game.writer.tracker.next_frame\[214\] net1336 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[214\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11691__A2 _05194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout168_A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13125__S net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11434__A game.CPU.applesa.ab.check_walls.above.walls\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_278_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09303_ net1085 game.CPU.applesa.ab.absxs.body_x\[55\] vssd1 vssd1 vccd1 vccd1 _03546_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_354_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout335_A game.CPU.walls.rand_wall.abduyd.next_wall\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16663__C _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1077_A game.CPU.applesa.x\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ game.CPU.applesa.ab.check_walls.above.walls\[190\] vssd1 vssd1 vccd1 vccd1
+ _03483_ sky130_fd_sc_hd__inv_2
XANTENNA__14464__B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10992__B net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_302_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12928__C1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09165_ game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1 vccd1 vccd1
+ _03414_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15590__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout123_X net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout502_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09096_ game.CPU.applesa.ab.absxs.body_y\[35\] vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_309_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_275_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09574__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_231_Right_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout871_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout969_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17095__B1 _02700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18924__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09293__B game.CPU.applesa.ab.check_walls.above.walls\[82\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09998_ game.CPU.apple_location\[1\] net1450 _04207_ vssd1 vssd1 vccd1 vccd1 _01366_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_71_Left_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14448__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08949_ net1129 vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_68_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__09324__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13751__S0 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09324__B2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ net573 _05198_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_240_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ net1166 _04808_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout924_X net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ net751 _05350_ _05355_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_357_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13630_ net247 _07503_ vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__nand2_1
XFILLER_0_211_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10842_ game.CPU.randy.counter1.count\[3\] _03513_ game.CPU.randy.counter1.count\[2\]
+ _03515_ _04744_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__o221a_1
XFILLER_0_183_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11063__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13561_ net201 _07426_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__or2_1
X_10773_ game.CPU.applesa.ab.absxs.body_y\[67\] _04679_ _04680_ net1270 vssd1 vssd1
+ vccd1 vccd1 _01014_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12631__B2 game.CPU.applesa.twoapples.absxs.next_head\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15300_ _08848_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12512_ game.CPU.applesa.ab.absxs.body_y\[74\] net522 net360 game.CPU.applesa.ab.absxs.body_y\[72\]
+ _06386_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__a221o_1
X_16280_ net872 _01516_ _02282_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__a21boi_2
X_13492_ _07105_ _07106_ _07116_ _07107_ net700 net489 vssd1 vssd1 vccd1 vccd1 _07366_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__14374__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17570__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15231_ game.CPU.applesa.normal1.number\[2\] _08790_ vssd1 vssd1 vccd1 vccd1 _08795_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_97_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17966__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12443_ game.CPU.applesa.ab.absxs.body_y\[107\] net366 net378 game.CPU.applesa.ab.absxs.body_x\[105\]
+ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_124_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12395__B1 game.CPU.applesa.twoapples.absxs.next_head\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_251_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15162_ net1213 net1239 game.CPU.applesa.ab.check_walls.above.walls\[190\] vssd1
+ vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__and3_1
X_12374_ _06247_ _06248_ _06249_ _06250_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__or4_1
XANTENNA__16125__A2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_300_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14113_ net882 game.CPU.applesa.ab.check_walls.above.walls\[169\] _03471_ net1052
+ vssd1 vssd1 vccd1 vccd1 _07987_ sky130_fd_sc_hd__o22a_1
XANTENNA__14136__A1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14136__B2 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325_ net815 net316 vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__and2_1
X_19970_ clknet_leaf_41_clk game.writer.tracker.next_frame\[565\] net1326 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[565\] sky130_fd_sc_hd__dfrtp_1
X_15093_ net1203 net1229 game.CPU.applesa.ab.check_walls.above.walls\[121\] vssd1
+ vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__and3_1
XANTENNA__12147__B1 _06026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14044_ net965 net943 vssd1 vssd1 vccd1 vccd1 _07918_ sky130_fd_sc_hd__or2_1
X_11256_ _05130_ _05143_ _05144_ _05145_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__or4b_4
X_18921_ clknet_leaf_5_clk net1390 _00605_ vssd1 vssd1 vccd1 vccd1 game.CPU.down_button.eD1.D
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17086__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _04392_ _04399_ _04393_ _04390_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__o211a_1
X_11187_ _03231_ net408 vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__xnor2_1
X_18852_ clknet_leaf_8_clk _01243_ _00562_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_274_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16833__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_340_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17803_ net870 _01566_ _03134_ _06633_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__o211a_1
XANTENNA__15492__Y _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ game.CPU.randy.f1.a1.count\[6\] game.CPU.randy.f1.a1.count\[4\] vssd1 vssd1
+ vccd1 vccd1 _04333_ sky130_fd_sc_hd__nand2_1
XANTENNA__11238__B net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15933__B net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18783_ clknet_leaf_10_clk _01200_ _00520_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[101\]
+ sky130_fd_sc_hd__dfrtp_1
X_15995_ game.CPU.applesa.ab.check_walls.above.walls\[97\] net472 net461 game.CPU.applesa.ab.check_walls.above.walls\[99\]
+ _02006_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_59_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
X_17734_ game.CPU.applesa.ab.count\[0\] net1167 vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__and2_1
X_10069_ _04240_ _04273_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__xnor2_1
X_14946_ _08719_ _08721_ _08722_ vssd1 vssd1 vccd1 vccd1 _08723_ sky130_fd_sc_hd__or3_1
XFILLER_0_221_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17665_ game.CPU.kyle.L1.cnt_500hz\[12\] _03053_ vssd1 vssd1 vccd1 vccd1 _03056_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_221_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14877_ game.CPU.walls.abc.number\[1\] game.CPU.walls.abc.number\[5\] game.CPU.walls.abc.counter
+ vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16616_ net156 _02370_ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__or2_1
X_19404_ clknet_leaf_70_clk _01404_ _00973_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.count1
+ sky130_fd_sc_hd__dfrtp_1
X_13828_ game.writer.tracker.frame\[539\] net708 net671 game.writer.tracker.frame\[540\]
+ _07701_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__o221a_1
X_17596_ _03002_ _03013_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16547_ net203 net146 _02396_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__and3_1
X_19335_ clknet_leaf_72_clk _01351_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.count_luck\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12784__S net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13759_ game.writer.tracker.frame\[131\] net708 net671 game.writer.tracker.frame\[132\]
+ vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_102_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19266_ clknet_leaf_8_clk _00054_ _00896_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_351_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16478_ net1702 _02426_ _02428_ _02273_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[60\]
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_333_Right_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18217_ net666 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__inv_2
XFILLER_0_289_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15429_ _01440_ _01455_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19197_ clknet_leaf_66_clk _00289_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.good_spot
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_31_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12085__A game.CPU.applesa.ab.check_walls.above.walls\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15099__C game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_215_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18148_ net627 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__inv_2
XANTENNA__17313__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_3_clk_X clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold203 game.writer.tracker.frame\[519\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 game.writer.tracker.frame\[293\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14127__A1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14127__B2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18947__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold225 game.writer.tracker.frame\[406\] vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_257_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18079_ net669 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__inv_2
Xhold236 game.writer.tracker.frame\[182\] vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 game.writer.tracker.frame\[184\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold258 game.writer.tracker.frame\[105\] vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 game.writer.tracker.frame\[409\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ net1262 _04152_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__nand2_1
XANTENNA__12689__A1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout705 net706 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__buf_4
XANTENNA__13886__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16004__B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout716 net717 vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__clkbuf_2
X_20041_ net1365 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__11429__A game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout727 net738 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_4
X_09852_ net1105 game.CPU.applesa.ab.absxs.body_x\[28\] vssd1 vssd1 vccd1 vccd1 _04095_
+ sky130_fd_sc_hd__nand2_1
Xfanout738 _04738_ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_4
XANTENNA__10333__A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_272_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout749 _04442_ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_237_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11148__B net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17092__A3 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_304_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ net910 game.CPU.applesa.ab.check_walls.above.walls\[144\] _03458_ net1154
+ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__a22o_1
XANTENNA__15843__B net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10620__X _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_252_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10987__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19104__Q game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout452_A net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1194_A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16674__B _02441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout240_X net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout717_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19722__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_315_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_300_Right_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14194__B net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09217_ game.CPU.applesa.ab.check_walls.above.walls\[162\] vssd1 vssd1 vccd1 vccd1
+ _03466_ sky130_fd_sc_hd__inv_2
XANTENNA__11611__B net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_279_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12377__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1247_X net1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09148_ game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1 vssd1 vccd1 vccd1
+ _03397_ sky130_fd_sc_hd__inv_2
XANTENNA__19930__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10388__C1 net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16107__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_295_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14118__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14118__B2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ game.CPU.applesa.ab.absxs.body_y\[83\] vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__inv_2
XANTENNA__16658__A3 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19872__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__A1_N net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11110_ _03347_ net533 vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_188_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12090_ _05973_ _05974_ _05975_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11041_ _03328_ game.CPU.applesa.ab.absxs.next_head\[7\] vssd1 vssd1 vccd1 vccd1
+ _04931_ sky130_fd_sc_hd__nor2_1
XANTENNA__11339__A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_338_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15753__B game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_271_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14800_ game.CPU.randy.counter1.count\[8\] _08612_ vssd1 vssd1 vccd1 vccd1 _08614_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_271_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _01788_ _01789_ _01790_ _01791_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__or4_1
XFILLER_0_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12992_ game.writer.tracker.frame\[574\] game.writer.tracker.frame\[575\] net1021
+ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09848__A2 game.CPU.applesa.ab.absxs.body_x\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14369__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14731_ game.CPU.randy.counter1.count1\[9\] _08559_ vssd1 vssd1 vccd1 vccd1 _08562_
+ sky130_fd_sc_hd__or2_1
X_11943_ net796 net310 vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__nand2_1
XANTENNA__11655__A2 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17240__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17450_ net612 _02879_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__nor2_1
X_14662_ game.CPU.randy.f1.state\[5\] game.CPU.randy.f1.state\[4\] _04345_ _08489_
+ vssd1 vssd1 vccd1 vccd1 _08501_ sky130_fd_sc_hd__o31a_1
X_11874_ game.CPU.applesa.ab.check_walls.above.walls\[140\] net390 vssd1 vssd1 vccd1
+ vccd1 _05762_ sky130_fd_sc_hd__nand2_1
X_16401_ net195 _02330_ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__nor2_4
X_13613_ net200 _07486_ net282 vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ _04482_ _04568_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nor2_1
X_17381_ _02787_ _02808_ _02810_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_253_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14593_ game.CPU.clock1.counter\[1\] game.CPU.clock1.counter\[0\] _08453_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.next_counter\[1\] sky130_fd_sc_hd__o21a_1
XANTENNA__13801__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19120_ net1182 _00160_ _00791_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[165\]
+ sky130_fd_sc_hd__dfrtp_4
X_16332_ net1986 net732 _02323_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[19\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__11802__A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13544_ net226 _07404_ net283 vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10756_ _04173_ _04593_ net329 vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_175_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19051_ net1191 _00283_ _00722_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[96\]
+ sky130_fd_sc_hd__dfrtp_2
X_16263_ _02230_ _02268_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__nor2_1
XANTENNA__11521__B net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13475_ net496 _07346_ _07348_ net214 vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__o211a_1
XFILLER_0_299_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16897__A3 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_341_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10687_ game.CPU.applesa.ab.absxs.body_y\[102\] _04595_ _04708_ game.CPU.applesa.ab.absxs.body_y\[98\]
+ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__a22o_1
X_18002_ net634 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__inv_2
X_15214_ game.CPU.applesa.normal1.number\[7\] _08775_ net758 vssd1 vssd1 vccd1 vccd1
+ _08781_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15487__Y net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12426_ game.CPU.applesa.ab.absxs.body_y\[102\] net519 vssd1 vssd1 vccd1 vccd1 _06303_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__19671__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15928__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16194_ _01823_ _01827_ _02060_ _02188_ _02205_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__o2111a_1
XANTENNA__10379__C1 net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09784__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15145_ net1216 net1236 game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1
+ vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__and3_1
XANTENNA__19600__RESET_B net1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16649__A3 _02413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12357_ game.CPU.applesa.ab.absxs.body_x\[45\] net379 vssd1 vssd1 vccd1 vccd1 _06234_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__09784__B2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ game.CPU.applesa.ab.check_walls.above.walls\[66\] net768 vssd1 vssd1 vccd1
+ vccd1 _05197_ sky130_fd_sc_hd__xor2_2
X_19953_ clknet_leaf_43_clk game.writer.tracker.next_frame\[548\] net1306 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[548\] sky130_fd_sc_hd__dfrtp_1
X_15076_ net1211 net1237 game.CPU.applesa.ab.check_walls.above.walls\[104\] vssd1
+ vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__and3_1
X_12288_ net830 net549 vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_264_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12352__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13332__A2 _06924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14027_ net877 game.CPU.applesa.ab.check_walls.above.walls\[162\] _07897_ _07898_
+ _07900_ vssd1 vssd1 vccd1 vccd1 _07901_ sky130_fd_sc_hd__a2111o_1
XANTENNA__09536__B2 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18904_ clknet_leaf_4_clk _01271_ _00588_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[2\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11249__A game.CPU.applesa.ab.absxs.body_y\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ game.CPU.applesa.ab.absxs.body_y\[111\] net398 vssd1 vssd1 vccd1 vccd1 _05129_
+ sky130_fd_sc_hd__nor2_1
X_19884_ clknet_leaf_26_clk game.writer.tracker.next_frame\[479\] net1312 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[479\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_248_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_206_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12540__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18835_ clknet_leaf_0_clk _01226_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18766_ clknet_leaf_51_clk _01183_ _00503_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[68\]
+ sky130_fd_sc_hd__dfrtp_4
X_15978_ game.CPU.applesa.ab.check_walls.above.walls\[68\] net453 vssd1 vssd1 vccd1
+ vccd1 _01990_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09839__A2 game.CPU.applesa.ab.absxs.body_y\[106\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_222_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17717_ net1998 _03086_ _03088_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__a21oi_1
X_14929_ _08705_ vssd1 vssd1 vccd1 vccd1 _08706_ sky130_fd_sc_hd__inv_2
XANTENNA__18553__RESET_B net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18697_ clknet_leaf_59_clk _01114_ _00434_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[43\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_353_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17648_ _03044_ _03037_ _03043_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__and3b_1
XANTENNA__19745__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_275_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17579_ net1437 net264 _03000_ _08809_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11712__A game.CPU.applesa.ab.apple_possible\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10606__B1 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09389__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19318_ clknet_leaf_71_clk _01342_ _00924_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.apple_location2_n\[2\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__16337__A2 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12527__B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_317_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11431__B net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19249_ clknet_leaf_7_clk _00063_ _00887_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__19895__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09002_ game.CPU.applesa.ab.absxs.body_x\[13\] vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_289_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13020__A1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_277_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15936__A1_N game.CPU.applesa.ab.check_walls.above.walls\[123\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15838__B net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_189_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10047__B net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13198__X _07072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__B2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout200_A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19125__CLK net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13308__C1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15848__A1 game.CPU.applesa.ab.absxs.body_x\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_286_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13859__B1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12262__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_284_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout502 net503 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_228_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09904_ _04120_ _04146_ net1079 net1263 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11159__A net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout513 net514 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__buf_2
XANTENNA__12757__S1 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16302__X _02301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12830__X _06704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout524 net527 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_4
XFILLER_0_272_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18230__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12531__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout535 net537 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_4
Xfanout546 _04814_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_6
XANTENNA__09852__A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20024_ net1277 vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
Xfanout557 net560 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__clkbuf_8
X_09835_ net917 game.CPU.applesa.ab.absxs.body_x\[105\] _03255_ net1111 _04077_ vssd1
+ vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__o221a_1
XANTENNA_input5_A gpio_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout568 _04460_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_308_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout190_X net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout579 net591 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_4
XANTENNA__19275__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10998__A game.CPU.applesa.ab.absxs.body_x\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16273__B2 _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ net910 game.CPU.applesa.ab.check_walls.above.walls\[96\] game.CPU.applesa.ab.check_walls.above.walls\[99\]
+ net924 _04006_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__a221o_1
XFILLER_0_308_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14189__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11606__B net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout834_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09697_ _03932_ _03933_ _03934_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__a211o_1
XFILLER_0_324_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09998__S _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_317_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14036__B1 game.CPU.applesa.ab.check_walls.above.walls\[115\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14587__A1 net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18673__Q game.CPU.applesa.ab.absxs.body_y\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_355_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_327_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12277__X _06163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11622__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610_ game.CPU.applesa.ab.absxs.body_x\[81\] _04673_ _04674_ game.CPU.applesa.ab.absxs.body_x\[77\]
+ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11590_ net743 _05478_ _05476_ net564 vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12437__B net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_308_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_289_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10541_ game.CPU.applesa.ab.absxs.body_x\[39\] _04642_ _04643_ game.CPU.applesa.ab.absxs.body_x\[35\]
+ vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__a22o_1
XANTENNA__14492__X _08366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13260_ _07130_ _07131_ _07132_ _07133_ net487 net682 vssd1 vssd1 vccd1 vccd1 _07134_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__15748__B net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10472_ _04602_ game.CPU.applesa.ab.absxs.body_x\[95\] _04601_ vssd1 vssd1 vccd1
+ vccd1 _01198_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12211_ _06005_ _06096_ _06007_ _06006_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__or4bb_1
XANTENNA__09766__A1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09766__B2 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13191_ net216 _07064_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_328_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12453__A game.CPU.applesa.ab.absxs.body_y\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12142_ net782 net552 vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__or2_1
XFILLER_0_349_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19618__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16950_ net163 _02396_ net88 _02656_ net1567 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[304\]
+ sky130_fd_sc_hd__a32o_1
X_12073_ net810 net551 vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__xor2_1
XANTENNA__16212__X _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ game.CPU.applesa.ab.absxs.body_x\[90\] net411 vssd1 vssd1 vccd1 vccd1 _04914_
+ sky130_fd_sc_hd__xnor2_1
X_15901_ game.CPU.applesa.ab.absxs.body_x\[42\] net469 vssd1 vssd1 vccd1 vccd1 _01913_
+ sky130_fd_sc_hd__xnor2_1
X_16881_ net178 net134 vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__nor2_1
XFILLER_0_218_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_244_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18620_ clknet_leaf_13_clk _01037_ _00357_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[114\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_216_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15832_ game.CPU.applesa.ab.absxs.body_y\[111\] net435 vssd1 vssd1 vccd1 vccd1 _01844_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__16803__A3 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14275__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18642__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19768__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18551_ clknet_leaf_45_clk _00974_ net1298 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.cmd_num\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_15763_ game.CPU.applesa.ab.absxs.body_y\[118\] net441 vssd1 vssd1 vccd1 vccd1 _01775_
+ sky130_fd_sc_hd__xnor2_1
X_12975_ _06640_ _06642_ net686 vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_339_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_234_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17502_ _02836_ _02857_ _02929_ _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__or4_1
X_14714_ _08549_ _08550_ net54 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__o21a_1
X_11926_ net748 _05507_ _05508_ net572 vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__a22o_1
X_18482_ net638 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__inv_2
X_15694_ game.CPU.applesa.ab.absxs.body_x\[30\] net465 vssd1 vssd1 vccd1 vccd1 _01706_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_358_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_346_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_234_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17433_ _02774_ net426 _02840_ _02838_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_123_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14645_ net1510 _08484_ _08485_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[21\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__15775__B1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11857_ net573 _05489_ _05490_ net751 vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__o22a_1
XANTENNA__18792__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12589__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15004__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13786__C1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17364_ net1116 _02792_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__or2_1
X_10808_ game.CPU.applesa.ab.absxs.body_y\[17\] _04699_ _04700_ game.CPU.applesa.ab.absxs.body_y\[13\]
+ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__a22o_1
XANTENNA__09454__B1 game.CPU.applesa.ab.absxs.body_y\[69\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14576_ game.CPU.clock1.counter\[11\] game.CPU.clock1.counter\[12\] game.CPU.clock1.counter\[18\]
+ game.CPU.clock1.counter\[10\] vssd1 vssd1 vccd1 vccd1 _08438_ sky130_fd_sc_hd__or4bb_1
X_11788_ net750 _05255_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__xnor2_1
X_16315_ _02244_ net236 net198 net203 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__and4b_4
XANTENNA__15498__X net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09002__A game.CPU.applesa.ab.absxs.body_x\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_184_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19103_ net1180 _00141_ _00774_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[148\]
+ sky130_fd_sc_hd__dfrtp_1
X_13527_ net995 net865 vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__nand2_2
X_17295_ net1919 net722 _02755_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[550\]
+ sky130_fd_sc_hd__and3_1
X_10739_ game.CPU.applesa.ab.absxs.body_y\[12\] _04653_ _04654_ game.CPU.applesa.ab.absxs.body_y\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11800__A2 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18315__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19034_ net1189 _00264_ _00705_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_16246_ _02228_ _02253_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__nor2_4
XFILLER_0_125_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ _06985_ _07017_ net704 vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__mux2_1
XANTENNA__15658__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_180_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_212_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11013__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ _03307_ net369 net521 game.CPU.applesa.ab.absxs.body_y\[54\] vssd1 vssd1
+ vccd1 vccd1 _06286_ sky130_fd_sc_hd__o22a_1
X_16177_ _03478_ net336 net439 game.CPU.applesa.ab.check_walls.above.walls\[182\]
+ _02027_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a221o_1
X_13389_ _07261_ _07262_ net481 vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10367__A2 _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15128_ net1208 net1233 game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1
+ vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__and3_1
XFILLER_0_266_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_259_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19298__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_254_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15674__A game.CPU.applesa.ab.check_walls.above.walls\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_19936_ clknet_leaf_42_clk game.writer.tracker.next_frame\[531\] net1326 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[531\] sky130_fd_sc_hd__dfrtp_1
X_15059_ net1211 net1242 net808 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__and3_1
XFILLER_0_254_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18050__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11316__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16489__B net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17047__A3 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19867_ clknet_leaf_20_clk game.writer.tracker.next_frame\[462\] net1308 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[462\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13906__B game.CPU.applesa.ab.check_walls.above.walls\[120\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09620_ net894 net832 net831 net908 _03862_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__a221o_1
XANTENNA__11707__A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_301_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18818_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[21\] _00555_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[21\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09391__B net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19798_ clknet_leaf_38_clk game.writer.tracker.next_frame\[393\] net1328 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[393\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_179_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_250_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_223_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09551_ net1111 _03256_ _03323_ net1149 _03793_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__a221o_1
XANTENNA__11426__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12816__A1 game.writer.tracker.frame\[329\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18749_ clknet_leaf_64_clk _01166_ _00486_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_222_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17204__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09482_ net915 game.CPU.applesa.ab.check_walls.above.walls\[177\] net783 net907 vssd1
+ vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_53_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout150_A net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13133__S net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_195_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12257__B net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_317_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_351_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_312_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout415_A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18225__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09847__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16191__B1 _01793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14472__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09566__B game.CPU.applesa.ab.absxs.body_y\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout203_X net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17286__A3 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09285__C _03527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout784_A game.CPU.applesa.ab.check_walls.above.walls\[180\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16032__X _02044_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1308 net1314 vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__clkbuf_4
Xfanout310 net311 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1112_X net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1319 net1323 vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__clkbuf_4
XANTENNA__18665__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout321 net323 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_4
Xfanout332 game.CPU.walls.rand_wall.abduyd.next_wall\[6\] vssd1 vssd1 vccd1 vccd1
+ net332 sky130_fd_sc_hd__buf_6
Xfanout343 game.CPU.walls.rand_wall.abduyd.next_wall\[3\] vssd1 vssd1 vccd1 vccd1
+ net343 sky130_fd_sc_hd__buf_6
XANTENNA__19910__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17038__A3 _02619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout354 net357 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout572_X net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout951_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_323_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12720__B net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout365 net366 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__buf_2
X_20007_ net1376 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
Xfanout376 _06209_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_2
Xfanout387 net389 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_4
X_09818_ net921 game.CPU.applesa.ab.absxs.body_x\[26\] _03348_ net1128 _04060_ vssd1
+ vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__a221o_1
XANTENNA__09920__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout398 net400 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14257__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout63_A net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10530__A2 _04609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09749_ _03983_ _03984_ _03988_ _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__or4_1
XANTENNA__11336__B net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_186_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12760_ net1065 _06551_ _06564_ _06579_ _06585_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__a32o_1
XFILLER_0_185_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14009__B1 game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17746__A1 game.CPU.applesa.ab.good_collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_328_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_295_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12719__Y _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11711_ net571 _04780_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__nand2_1
XANTENNA__17023__B _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17210__A3 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12691_ _06561_ _06563_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__xor2_4
XANTENNA__13043__S net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14430_ _08301_ _08303_ vssd1 vssd1 vccd1 vccd1 _08304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ game.CPU.applesa.ab.check_walls.above.walls\[158\] net254 vssd1 vssd1 vccd1
+ vccd1 _05531_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_327_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_315_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16862__B _02415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12167__B net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15759__A game.CPU.applesa.ab.absxs.body_y\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14361_ game.CPU.applesa.ab.absxs.body_x\[101\] net884 net1055 _03227_ vssd1 vssd1
+ vccd1 vccd1 _08235_ sky130_fd_sc_hd__a22o_1
X_11573_ net773 _05461_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16100_ _01839_ _01840_ _02110_ _02111_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__or4b_1
X_13312_ _06744_ _06753_ _06755_ _06754_ net505 net696 vssd1 vssd1 vccd1 vccd1 _07186_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17080_ _02467_ net57 _02696_ net1618 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[394\]
+ sky130_fd_sc_hd__a22o_1
X_10524_ net934 game.CPU.applesa.ab.absxs.body_x\[56\] vssd1 vssd1 vccd1 vccd1 _04636_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09757__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14292_ game.CPU.applesa.ab.absxs.body_y\[54\] net957 vssd1 vssd1 vccd1 vccd1 _08166_
+ sky130_fd_sc_hd__xor2_1
Xwire755 _03528_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14382__B net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16031_ _03296_ net333 vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13243_ game.writer.tracker.frame\[500\] game.writer.tracker.frame\[501\] net1014
+ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__mux2_1
XANTENNA__19440__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ net850 _04588_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__or2_4
X_13174_ game.writer.tracker.frame\[448\] game.writer.tracker.frame\[449\] net1039
+ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__mux2_2
X_10386_ net1153 game.CPU.apple_location\[4\] vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__and2_1
XFILLER_0_248_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_248_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16485__A1 _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_43_clk_X clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ _06009_ _06010_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__or3b_2
XFILLER_0_248_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12911__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_176_Right_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17982_ net606 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__inv_2
XFILLER_0_263_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_261_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19590__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19721_ clknet_leaf_24_clk game.writer.tracker.next_frame\[316\] net1346 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[316\] sky130_fd_sc_hd__dfrtp_1
X_16933_ net184 _02521_ net87 _02651_ net1537 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[292\]
+ sky130_fd_sc_hd__a32o_1
X_12056_ _05440_ _05441_ _05444_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__nor3_1
XANTENNA__16237__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16102__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _03308_ net536 vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15781__X _01793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11527__A net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19652_ clknet_leaf_21_clk game.writer.tracker.next_frame\[247\] net1343 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[247\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15450__D_N net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16864_ _02544_ net107 _02626_ net1852 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[247\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_125_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14248__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16788__A2 _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_58_clk_X clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_245_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18603_ clknet_leaf_3_clk _00005_ _00340_ vssd1 vssd1 vccd1 vccd1 game.CPU.luck1.Qa\[0\]
+ sky130_fd_sc_hd__dfstp_4
XANTENNA__15941__B net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15815_ _01824_ _01825_ _01826_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__or3_1
X_19583_ clknet_leaf_34_clk game.writer.tracker.next_frame\[178\] net1338 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[178\] sky130_fd_sc_hd__dfrtp_1
X_16795_ _02475_ net102 _02599_ net1526 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[206\]
+ sky130_fd_sc_hd__a22o_1
X_15746_ game.CPU.applesa.ab.check_walls.above.walls\[1\] net473 vssd1 vssd1 vccd1
+ vccd1 _01758_ sky130_fd_sc_hd__xnor2_1
X_18534_ net628 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__inv_2
X_12958_ net224 _06756_ _06831_ net274 vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_319_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_259_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11909_ net573 _05282_ _05286_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_358_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17201__A3 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15677_ game.CPU.applesa.ab.check_walls.above.walls\[15\] net434 vssd1 vssd1 vccd1
+ vccd1 _01689_ sky130_fd_sc_hd__xor2_1
X_18465_ net652 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12889_ game.writer.tracker.frame\[60\] game.writer.tracker.frame\[61\] net1040 vssd1
+ vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__mux2_1
XANTENNA__12358__A game.CPU.applesa.ab.absxs.body_x\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_272_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14628_ game.CPU.clock1.counter\[15\] _08474_ vssd1 vssd1 vccd1 vccd1 _08475_ sky130_fd_sc_hd__and2_1
X_17416_ _08443_ _02778_ net426 vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__and3b_1
XFILLER_0_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18396_ net617 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10037__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17347_ _02771_ _02776_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__nand2_1
XANTENNA__13774__A2 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14971__A1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14559_ net1176 game.CPU.walls.abc.number_out\[5\] vssd1 vssd1 vccd1 vccd1 _08426_
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_333_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14971__B2 net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12645__X _06522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10588__A2 _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_302_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09667__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17278_ net176 _02258_ _02341_ _02750_ net1795 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[538\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_12_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16173__B1 game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16712__A2 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14292__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_348_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16229_ net175 net132 vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__nor2_4
X_19017_ net1193 _00246_ _00688_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[62\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12734__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19933__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_283_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08982_ game.CPU.applesa.ab.absxs.body_x\[87\] vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__inv_2
XFILLER_0_255_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_225_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_299_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19919_ clknet_leaf_33_clk game.writer.tracker.next_frame\[514\] net1301 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[514\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_254_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16012__B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout198_A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13128__S net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__A1 _03677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16779__A2 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ _03837_ _03838_ _03844_ _03845_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__a22o_1
XANTENNA__11156__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15851__B net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ game.CPU.applesa.ab.snake_head_x\[2\] game.CPU.applesa.ab.check_walls.above.walls\[74\]
+ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__xor2_1
XFILLER_0_167_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10995__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_210_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09465_ net1098 game.CPU.applesa.ab.absxs.body_x\[93\] vssd1 vssd1 vccd1 vccd1 _03708_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__19112__Q game.CPU.applesa.ab.check_walls.above.walls\[157\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09396_ net1084 game.CPU.applesa.ab.check_walls.above.walls\[91\] vssd1 vssd1 vccd1
+ vccd1 _03639_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14411__B1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13765__A2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1062_X net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_278_Right_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10579__A2 game.CPU.applesa.ab.absxs.body_x\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09577__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13099__A net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_332_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17794__A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__S0 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11528__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1327_X net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10240_ _04377_ _04429_ _04403_ _04380_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_325_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17259__A3 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ _04363_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_245_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14478__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10751__A2 _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1105 net1106 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_273_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1116 game.CPU.bodymain1.main.score\[4\] vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__buf_2
Xfanout1127 net1129 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout954_X net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1138 game.CPU.applesa.ab.snake_head_y\[2\] vssd1 vssd1 vccd1 vccd1 net1138
+ sky130_fd_sc_hd__buf_4
Xfanout151 _02270_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_261_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12450__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1149 net1151 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__buf_4
Xfanout162 _06701_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_4
XANTENNA__13038__S net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13930_ net961 net823 vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__or2_1
Xfanout173 _06702_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_4
XANTENNA__10251__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout184 net187 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_346_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout195 net196 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_6
XANTENNA__09462__D net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10503__A2 _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13861_ net274 _07731_ _07734_ net506 vssd1 vssd1 vccd1 vccd1 _07735_ sky130_fd_sc_hd__a211o_1
XANTENNA__15761__B net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15600_ game.CPU.applesa.ab.check_walls.above.walls\[113\] net471 net343 _03441_
+ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__a22o_1
X_12812_ game.writer.tracker.frame\[362\] game.writer.tracker.frame\[363\] net1001
+ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__mux2_1
X_16580_ _02340_ _02493_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_18_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13792_ _07664_ _07665_ net484 vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_336_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14377__B net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15531_ _01531_ _01550_ _01552_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_70_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ _06615_ _06616_ net488 vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__mux2_1
XANTENNA__19444__RESET_B net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19806__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17195__A2 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19022__Q game.CPU.applesa.ab.check_walls.above.walls\[67\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18250_ net622 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
X_15462_ _01440_ _01450_ _01454_ _01462_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__or4_1
XFILLER_0_166_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12674_ game.writer.control.current\[0\] game.writer.control.current\[1\] vssd1 vssd1
+ vccd1 vccd1 _06548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17201_ net56 _02439_ net74 _02731_ net1598 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[480\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_181_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14413_ game.CPU.applesa.ab.absxs.body_x\[45\] net884 net854 game.CPU.applesa.ab.absxs.body_y\[46\]
+ vssd1 vssd1 vccd1 vccd1 _08287_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__15489__A _08368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11625_ game.CPU.applesa.ab.check_walls.above.walls\[190\] net254 vssd1 vssd1 vccd1
+ vccd1 _05514_ sky130_fd_sc_hd__xnor2_1
X_18181_ net609 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__inv_2
X_15393_ game.writer.updater.commands.mode\[2\] game.writer.updater.commands.mode\[1\]
+ game.writer.updater.commands.mode\[0\] vssd1 vssd1 vccd1 vccd1 _08935_ sky130_fd_sc_hd__or3b_2
XFILLER_0_181_132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12964__B1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17132_ _02310_ net165 net76 _02712_ net1601 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[430\]
+ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_245_Right_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_343_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09487__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14344_ _03244_ net1055 net869 game.CPU.applesa.ab.absxs.body_y\[36\] _08216_ vssd1
+ vssd1 vccd1 vccd1 _08218_ sky130_fd_sc_hd__a221o_1
X_11556_ _04460_ _05440_ _05441_ net743 vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__a22o_1
XANTENNA__18830__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19956__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11404__A1_N game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17063_ _02436_ net83 _02689_ net1558 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[384\]
+ sky130_fd_sc_hd__a22o_1
X_10507_ net754 _04606_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__nor2_4
X_14275_ game.CPU.applesa.ab.absxs.body_x\[48\] net889 net1056 _03272_ vssd1 vssd1
+ vccd1 vccd1 _08149_ sky130_fd_sc_hd__o22a_1
XANTENNA__15001__B net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11487_ game.CPU.applesa.ab.check_walls.above.walls\[54\] net256 _05372_ _05373_
+ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__o2111a_1
XANTENNA__11519__A1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16014_ game.CPU.applesa.ab.check_walls.above.walls\[176\] net357 vssd1 vssd1 vccd1
+ vccd1 _02026_ sky130_fd_sc_hd__xnor2_1
X_13226_ _07095_ _07098_ net690 vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10438_ net1449 net847 _04161_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__a21o_1
XANTENNA__14181__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18980__CLK net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ game.writer.tracker.frame\[156\] game.writer.tracker.frame\[157\] net1035
+ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09934__B _03527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10369_ game.CPU.applesa.ab.absxs.body_y\[4\] net847 _04158_ net1451 vssd1 vssd1
+ vccd1 vccd1 _01273_ sky130_fd_sc_hd__a22o_1
XFILLER_0_236_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12108_ net819 net290 vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__xor2_1
X_13088_ _06960_ _06961_ net477 vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__mux2_1
X_17965_ net668 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__inv_2
XFILLER_0_291_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12360__B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19704_ clknet_leaf_31_clk game.writer.tracker.next_frame\[299\] net1281 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[299\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15952__A game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16916_ net69 _02643_ _02647_ net1884 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[279\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12039_ net801 net289 vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__nor2_1
XFILLER_0_256_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_251_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09896__B1 _04138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19336__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17896_ net643 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__inv_2
XFILLER_0_217_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19635_ clknet_leaf_28_clk game.writer.tracker.next_frame\[230\] net1290 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[230\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15671__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16847_ net131 _02389_ net143 vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_252_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16630__A1 _02299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_220_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19566_ clknet_leaf_38_clk game.writer.tracker.next_frame\[161\] net1328 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[161\] sky130_fd_sc_hd__dfrtp_2
X_16778_ _02450_ net108 _02594_ net1762 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[194\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_38_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18517_ net581 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__inv_2
XANTENNA__11455__B1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19486__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15729_ _03319_ net337 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__xnor2_1
X_19497_ clknet_leaf_25_clk game.writer.tracker.next_frame\[92\] net1321 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[92\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12088__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17186__A2 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09250_ game.CPU.randy.counter1.count\[15\] vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__inv_2
X_18448_ net592 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__inv_2
XANTENNA__16933__A2 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18771__Q game.CPU.applesa.ab.absxs.body_x\[77\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13747__A2 game.writer.tracker.frame\[176\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_192_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09181_ net805 vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__inv_2
X_18379_ net600 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11758__B2 game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09397__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_212_Right_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload52_A clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16697__A1 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_231_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout113_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18503__A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13380__B1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12551__A game.CPU.applesa.ab.absxs.body_y\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17110__A2 _02434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1022_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_227_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11265__A2_N net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ net1206 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout482_A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12270__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15862__A game.CPU.applesa.ab.absxs.body_x\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_320_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09887__B1 _04129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15581__B net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_316_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout270_X net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19829__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18703__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_347_Right_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13435__A1 _06967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_316_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09517_ net1159 game.CPU.applesa.ab.absxs.body_y\[48\] vssd1 vssd1 vccd1 vccd1 _03760_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_39_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_292_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout914_A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout535_X net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11997__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_332_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11997__B2 game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ net914 game.CPU.applesa.ab.check_walls.above.walls\[137\] _03452_ net1089
+ _03690_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__o221a_1
XANTENNA__18853__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16924__A2 _02643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17301__B net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ net1131 net829 vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_156_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12726__A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_331_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12946__B1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11749__B2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ net797 net255 _05297_ _05298_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16137__B1 _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12390_ _03281_ game.CPU.applesa.twoapples.absxs.next_head\[0\] vssd1 vssd1 vccd1
+ vccd1 _06267_ sky130_fd_sc_hd__nor2_1
XANTENNA__12410__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10517__Y _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16688__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09100__A game.CPU.applesa.ab.absxs.body_y\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14148__C1 _08021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11341_ net564 _05224_ _05225_ _05229_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__o211a_1
X_14060_ net1060 game.CPU.applesa.ab.check_walls.above.walls\[145\] vssd1 vssd1 vccd1
+ vccd1 _07934_ sky130_fd_sc_hd__xor2_1
XFILLER_0_277_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15756__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11272_ _05154_ _05158_ _05161_ _04875_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__o211a_1
XFILLER_0_278_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12174__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_320_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13011_ game.writer.tracker.frame\[524\] game.writer.tracker.frame\[525\] net1004
+ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_320_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10223_ _04404_ _04414_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09754__B net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10533__X _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_245_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19359__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13349__S1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ game.CPU.randy.f1.state\[1\] game.CPU.randy.f1.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _04349_ sky130_fd_sc_hd__and2_1
XFILLER_0_357_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19017__Q game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16860__A1 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15772__A game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_206_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17750_ net1271 _04304_ _03107_ _03108_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__o211ai_4
X_14962_ _08711_ _08720_ _08709_ vssd1 vssd1 vccd1 vccd1 _08739_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_233_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10085_ _04214_ _04222_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__or2_1
Xhold7 game.CPU.left_button.eD1.D vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__dlygate4sd3_1
X_16701_ _02477_ net63 _02567_ game.writer.tracker.frame\[144\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[144\] sky130_fd_sc_hd__a22o_1
X_13913_ net1052 _03445_ game.CPU.applesa.ab.check_walls.above.walls\[124\] net867
+ vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14893_ net1096 _08417_ vssd1 vssd1 vccd1 vccd1 _08670_ sky130_fd_sc_hd__and2_1
X_17681_ game.CPU.walls.rand_wall.count_luck\[1\] _03063_ net1749 vssd1 vssd1 vccd1
+ vccd1 _03067_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_226_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19420_ clknet_leaf_48_clk game.writer.tracker.next_frame\[15\] net1303 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13844_ net481 _07714_ _07715_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__and3_1
X_16632_ net53 _02518_ _02534_ net1730 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[108\]
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_314_Right_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_348_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19351_ clknet_leaf_71_clk game.CPU.applesa.twoapples.absxs.next_head\[7\] vssd1
+ vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.y_final\[3\] sky130_fd_sc_hd__dfxtp_1
X_13775_ net498 _07647_ _07648_ net231 vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__a31o_1
X_16563_ net225 _02411_ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__nor2_4
XFILLER_0_97_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10987_ game.CPU.applesa.ab.absxs.body_y\[112\] net536 vssd1 vssd1 vccd1 vccd1 _04877_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_48_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_256_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18302_ net643 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
X_12726_ net841 net840 vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__nand2_2
X_15514_ _01470_ _01536_ _01522_ _01492_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11988__B2 game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16494_ net190 net171 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__nand2_1
X_19282_ clknet_leaf_67_clk _01331_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.count\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_242_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15445_ _08396_ _01471_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_178_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18233_ net649 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__inv_2
X_12657_ game.CPU.applesa.ab.absxs.body_x\[66\] net373 game.CPU.applesa.twoapples.absxs.next_head\[4\]
+ _03336_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__a22o_1
XANTENNA__10660__B2 game.CPU.applesa.ab.absxs.body_x\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11608_ net565 _05491_ _05496_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__a21o_1
XANTENNA__15012__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15376_ _08913_ _08917_ vssd1 vssd1 vccd1 vccd1 _08918_ sky130_fd_sc_hd__or2_1
XANTENNA__16128__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18164_ net633 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__inv_2
X_12588_ net1268 net528 net370 game.CPU.applesa.ab.absxs.body_x\[90\] vssd1 vssd1
+ vccd1 vccd1 _06465_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12355__B game.CPU.applesa.twoapples.absxs.next_head\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17115_ net1886 _02706_ _02707_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[418\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14327_ game.CPU.applesa.ab.absxs.body_y\[75\] net941 vssd1 vssd1 vccd1 vccd1 _08201_
+ sky130_fd_sc_hd__or2_1
X_11539_ _05427_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__inv_2
X_18095_ net606 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold407 game.writer.tracker.frame\[450\] vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold418 game.writer.tracker.frame\[255\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_345_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17046_ _02321_ _02678_ net557 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold429 game.writer.tracker.frame\[104\] vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
X_14258_ game.CPU.applesa.ab.absxs.body_y\[79\] net941 vssd1 vssd1 vccd1 vccd1 _08132_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_311_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13209_ game.writer.tracker.frame\[426\] game.writer.tracker.frame\[427\] net1020
+ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_267_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12371__A game.CPU.applesa.ab.absxs.body_x\[115\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14189_ game.CPU.applesa.ab.absxs.body_y\[98\] net949 vssd1 vssd1 vccd1 vccd1 _08063_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10715__A2 _04609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout909 _03199_ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11912__A1 game.CPU.applesa.ab.check_walls.above.walls\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_209_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11912__B2 game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18997_ net1194 _00224_ _00668_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[42\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__18726__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15682__A game.CPU.applesa.ab.absxs.body_y\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17948_ net639 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_0_Left_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09680__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17879_ net656 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16603__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11274__X _05164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19618_ clknet_leaf_22_clk game.writer.tracker.next_frame\[213\] net1337 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[213\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_283_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_356_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18876__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16784__Y _02597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11691__A3 _05206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19549_ clknet_leaf_34_clk game.writer.tracker.next_frame\[144\] net1328 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[144\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__11434__B net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_278_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09302_ _03539_ _03542_ _03543_ _03544_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13930__A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12640__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ game.CPU.applesa.ab.check_walls.above.walls\[189\] vssd1 vssd1 vccd1 vccd1
+ _03482_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10651__A1 game.CPU.applesa.ab.absxs.body_x\[40\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout230_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_307_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11450__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16119__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09164_ net817 vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__inv_2
XFILLER_0_302_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12265__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15590__B2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09095_ game.CPU.applesa.ab.absxs.body_y\[40\] vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__inv_2
XFILLER_0_287_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18233__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_287_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1237_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19501__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09855__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_309_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15576__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_287_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout697_A net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12281__A game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1025_X net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10706__A2 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17095__A1 _02489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ game.CPU.apple_location\[2\] game.CPU.applesa.ab.apple_location\[2\] _04207_
+ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_A net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19651__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ net1119 vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__inv_2
XFILLER_0_215_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18676__Q game.CPU.applesa.ab.absxs.body_x\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_215_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_240_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ net1271 game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nor2_4
XANTENNA__13408__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_230_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11890_ _03389_ net309 vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_343_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10841_ game.CPU.randy.counter1.count\[2\] _03515_ game.CPU.randy.counter1.count\[1\]
+ _03517_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_333_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ net476 _07432_ _07433_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__and3_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ game.CPU.applesa.ab.absxs.body_y\[72\] _04675_ _04676_ game.CPU.applesa.ab.absxs.body_y\[68\]
+ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__a22o_1
X_12511_ game.CPU.applesa.ab.absxs.body_x\[75\] net531 game.CPU.applesa.twoapples.absxs.next_head\[4\]
+ _03333_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__a22o_1
XANTENNA__14908__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10642__A1 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13491_ net487 _07153_ _07364_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12919__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15230_ game.CPU.applesa.normal1.number\[6\] _08788_ vssd1 vssd1 vccd1 vccd1 _08794_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ _03252_ game.CPU.applesa.twoapples.absxs.next_head\[3\] game.CPU.applesa.twoapples.absxs.next_head\[4\]
+ _03321_ _06318_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_97_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_325_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13041__C1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_205_Left_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_288_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15161_ net1213 net1239 game.CPU.applesa.ab.check_walls.above.walls\[189\] vssd1
+ vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_251_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12373_ game.CPU.applesa.ab.absxs.body_x\[113\] net378 net361 game.CPU.applesa.ab.absxs.body_y\[112\]
+ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08940__Y _03190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14112_ net1062 _03470_ _03472_ net1043 vssd1 vssd1 vccd1 vccd1 _07986_ sky130_fd_sc_hd__o22a_1
XANTENNA__19181__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11324_ net563 _05192_ _05212_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__o21a_2
XANTENNA__09765__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15092_ net1203 net1229 game.CPU.applesa.ab.check_walls.above.walls\[120\] vssd1
+ vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18749__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14043_ net993 net954 vssd1 vssd1 vccd1 vccd1 _07917_ sky130_fd_sc_hd__nor2_1
X_18920_ clknet_leaf_5_clk net6 _00604_ vssd1 vssd1 vccd1 vccd1 game.CPU.down_button.sync1.Q
+ sky130_fd_sc_hd__dfrtp_1
X_11255_ game.CPU.applesa.ab.absxs.body_x\[111\] net546 net539 game.CPU.applesa.ab.absxs.body_y\[110\]
+ _05134_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__o221a_1
XANTENNA__12191__A game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19877__RESET_B net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13895__A1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17086__A1 _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13895__B2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ _04390_ _04395_ _04398_ _04397_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__a31oi_2
X_18851_ clknet_leaf_8_clk _01242_ _00561_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_11186_ game.CPU.applesa.ab.absxs.body_y\[86\] net403 vssd1 vssd1 vccd1 vccd1 _05076_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_207_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16294__C1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17802_ net696 _03138_ _03139_ net966 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__a22o_1
X_10137_ _04326_ _04329_ _04330_ _04331_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_214_Left_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18782_ clknet_leaf_10_clk _01199_ _00519_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[100\]
+ sky130_fd_sc_hd__dfrtp_4
X_15994_ game.CPU.applesa.ab.check_walls.above.walls\[101\] net444 vssd1 vssd1 vccd1
+ vccd1 _02006_ sky130_fd_sc_hd__xnor2_1
X_17733_ _03085_ _03098_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__nor2_1
XANTENNA__11658__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18586__Q game.CPU.applesa.ab.absxs.body_y\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_206_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10068_ _04219_ _04222_ _04227_ _04275_ _04229_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__a221o_1
X_14945_ _08676_ _08683_ _08718_ vssd1 vssd1 vccd1 vccd1 _08722_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13226__S net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15007__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17664_ game.CPU.kyle.L1.cnt_500hz\[12\] _03053_ vssd1 vssd1 vccd1 vccd1 _03055_
+ sky130_fd_sc_hd__or2_1
X_14876_ game.CPU.walls.abc.number\[0\] game.CPU.walls.abc.number\[4\] game.CPU.walls.abc.counter
+ vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_253_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19403_ clknet_leaf_47_clk _01403_ net1280 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.x\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_16615_ _02522_ _02524_ _02523_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[101\]
+ sky130_fd_sc_hd__a21o_1
X_13827_ game.writer.tracker.frame\[538\] net845 net835 game.writer.tracker.frame\[537\]
+ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__o22a_1
X_17595_ game.CPU.kyle.L1.cnt_20ms\[3\] _03001_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__nor2_1
XANTENNA__11822__X _05710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19334_ clknet_leaf_71_clk _01350_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.count_luck\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_16546_ net207 _02396_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__and2_2
X_13758_ game.writer.tracker.frame\[134\] net841 net834 game.writer.tracker.frame\[133\]
+ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__o22a_1
XANTENNA__17546__C1 _00293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12709_ _06578_ _06582_ _06566_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10633__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19265_ clknet_leaf_8_clk _00053_ _00895_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_16477_ _02254_ _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__nor2_8
X_13689_ _07554_ _07555_ _07562_ net277 net246 vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_223_Left_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_351_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18216_ net664 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19524__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15428_ _01449_ _01454_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__or2_1
XANTENNA__14375__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13032__C1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19196_ clknet_leaf_46_clk game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1
+ vccd1 vccd1 game.CPU.walls.rand_wall.y_final\[3\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_289_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12085__B net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15359_ _03366_ _08881_ vssd1 vssd1 vccd1 vccd1 _08901_ sky130_fd_sc_hd__xnor2_1
X_18147_ net626 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_215_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14581__A net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold204 game.writer.tracker.frame\[343\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09675__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold215 game.writer.tracker.frame\[282\] vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold226 game.writer.tracker.frame\[146\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ net669 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__inv_2
Xhold237 game.writer.tracker.frame\[116\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__A1 game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_348_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19674__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold248 game.CPU.applesa.apple_location2_n\[6\] vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15875__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12138__B2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09920_ net1084 net847 _04161_ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__a21o_1
X_17029_ net68 _02678_ _02680_ net1587 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[359\]
+ sky130_fd_sc_hd__a22o_1
Xhold259 game.CPU.randy.f1.a1.count\[5\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13886__A1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13886__B2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17077__A1 _02464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout706 net707 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_2
X_20040_ net1364 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout717 net726 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__clkbuf_4
X_09851_ net1105 game.CPU.applesa.ab.absxs.body_x\[28\] vssd1 vssd1 vccd1 vccd1 _04094_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_113_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout728 net738 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11429__B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_232_Left_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19547__RESET_B net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout739 _04486_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkload15_A clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09782_ net1145 game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1 vccd1
+ vccd1 _04025_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_304_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16020__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10872__A1 game.CPU.randy.counter1.count\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19054__CLK net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12975__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14063__A1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14063__B2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout445_A _08427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1187_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17001__A1 _02486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09490__A1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout612_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19120__Q game.CPU.applesa.ab.check_walls.above.walls\[165\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12276__A game.CPU.applesa.ab.check_walls.above.walls\[159\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_315_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09490__B2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11180__A game.CPU.applesa.ab.absxs.body_y\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09216_ game.CPU.applesa.ab.check_walls.above.walls\[161\] vssd1 vssd1 vccd1 vccd1
+ _03465_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_350_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09147_ game.CPU.applesa.ab.check_walls.above.walls\[32\] vssd1 vssd1 vccd1 vccd1
+ _03396_ sky130_fd_sc_hd__inv_2
XFILLER_0_322_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1142_X net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09585__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ game.CPU.applesa.ab.absxs.body_y\[88\] vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout981_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13877__A1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout93_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13877__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ _04923_ _04928_ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_34_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_235_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11888__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10560__B1 _04652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ game.writer.tracker.frame\[570\] game.writer.tracker.frame\[571\] net1021
+ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_271_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11355__A game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11942_ net787 net300 _05820_ _05821_ _05829_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__o2111a_1
X_14730_ game.CPU.randy.counter1.count1\[9\] _08559_ vssd1 vssd1 vccd1 vccd1 _08561_
+ sky130_fd_sc_hd__and2_1
XANTENNA__16579__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17240__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11074__B net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14661_ net752 _08499_ vssd1 vssd1 vccd1 vccd1 _08500_ sky130_fd_sc_hd__or2_1
X_11873_ game.CPU.applesa.ab.check_walls.above.walls\[140\] net390 vssd1 vssd1 vccd1
+ vccd1 _05761_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15251__B1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16400_ net199 net165 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__nand2_2
X_13612_ _07484_ _07485_ net500 vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10824_ net1274 net1273 _04733_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__mux2_1
X_14592_ game.CPU.clock1.counter\[1\] game.CPU.clock1.counter\[0\] net739 vssd1 vssd1
+ vccd1 vccd1 _08453_ sky130_fd_sc_hd__a21oi_1
X_17380_ _02801_ _02804_ _02809_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_45_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_253_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10615__A1 game.CPU.applesa.ab.absxs.body_x\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13543_ net492 _07407_ _07408_ _07409_ net212 vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__a311o_1
X_16331_ net1959 net732 _02323_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[18\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__11802__B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10755_ game.CPU.applesa.ab.absxs.body_y\[108\] _04665_ _04666_ game.CPU.applesa.ab.absxs.body_y\[104\]
+ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__a22o_1
XANTENNA__10258__X _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17977__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11812__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16881__A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09481__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09481__B2 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16262_ net183 _02228_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__nor2_1
X_19050_ net1185 _00282_ _00721_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[95\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13474_ net512 _07347_ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__or2_1
X_10686_ game.CPU.applesa.ab.absxs.body_y\[103\] _04595_ _04708_ game.CPU.applesa.ab.absxs.body_y\[99\]
+ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_299_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15213_ game.CPU.applesa.normal1.number\[7\] _08775_ vssd1 vssd1 vccd1 vccd1 _08780_
+ sky130_fd_sc_hd__or2_1
X_18001_ net614 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__inv_2
XFILLER_0_341_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19697__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12425_ _06292_ _06301_ _06294_ _06298_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__or4b_1
X_16193_ _01778_ _01781_ _02196_ _02204_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10918__A2 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_301_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15144_ net1210 net1235 net785 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__and3_1
XANTENNA__09495__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ game.CPU.applesa.ab.absxs.body_x\[77\] net377 vssd1 vssd1 vccd1 vccd1 _06233_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ game.CPU.applesa.ab.check_walls.above.walls\[71\] net260 vssd1 vssd1 vccd1
+ vccd1 _05196_ sky130_fd_sc_hd__xnor2_1
X_19952_ clknet_leaf_43_clk game.writer.tracker.next_frame\[547\] net1306 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[547\] sky130_fd_sc_hd__dfrtp_1
X_15075_ net1212 net1238 net802 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__and3_1
X_12287_ _06169_ _06170_ _06171_ _06172_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__or4_2
XFILLER_0_239_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17059__A1 _02429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_264_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14026_ net886 game.CPU.applesa.ab.check_walls.above.walls\[160\] game.CPU.applesa.ab.check_walls.above.walls\[163\]
+ net876 _07899_ vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__a221o_1
X_18903_ clknet_leaf_4_clk _01270_ _00587_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11238_ game.CPU.applesa.ab.absxs.body_y\[111\] net398 vssd1 vssd1 vccd1 vccd1 _05128_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11249__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19883_ clknet_leaf_26_clk game.writer.tracker.next_frame\[478\] net1312 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[478\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11879__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15944__B game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11343__A2 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18834_ clknet_leaf_0_clk _01225_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11169_ game.CPU.applesa.ab.absxs.body_y\[76\] net534 vssd1 vssd1 vccd1 vccd1 _05059_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18765_ clknet_leaf_51_clk _01182_ _00502_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[63\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__19077__CLK net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15977_ _01977_ _01978_ _01987_ _01988_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17716_ game.CPU.applesa.ab.count_luck\[1\] _03086_ _03085_ vssd1 vssd1 vccd1 vccd1
+ _03088_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_165_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14928_ _08660_ _08703_ _08663_ vssd1 vssd1 vccd1 vccd1 _08705_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_264_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18696_ clknet_leaf_59_clk _01113_ _00433_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[42\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17231__A1 _02544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_353_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_348_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_90_Left_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17647_ game.CPU.kyle.L1.cnt_500hz\[6\] _08804_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__and2_1
X_14859_ _08649_ _08650_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[12\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_348_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13480__A net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_275_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17578_ _02772_ _02778_ _02827_ _02872_ _02878_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__a311oi_1
XANTENNA__16990__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19317_ clknet_leaf_71_clk _01341_ _00923_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.apple_location2_n\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_16529_ net149 net125 _02466_ _02463_ net2013 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[73\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17887__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09389__B game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09472__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18914__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09472__B2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16337__A3 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17534__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_332_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_317_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19248_ clknet_leaf_17_clk _00062_ _00886_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09001_ game.CPU.applesa.ab.absxs.body_x\[21\] vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__inv_2
XANTENNA__13556__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19179_ clknet_leaf_6_clk _01298_ _00841_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_189_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09775__A2 game.CPU.applesa.ab.YMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19728__RESET_B net1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_285_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16015__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12543__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15848__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_257_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_286_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18511__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09903_ _04128_ _04137_ _04141_ _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__and4_1
XFILLER_0_245_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout503 net516 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_228_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15854__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11159__B net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout514 net515 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout525 net527 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout536 net537 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_272_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09834_ net1149 game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1 vccd1 vccd1 _04077_
+ sky130_fd_sc_hd__xnor2_1
Xfanout547 net548 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_4
X_20023_ net1277 vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09852__B game.CPU.applesa.ab.absxs.body_x\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout558 net559 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1102_A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 net570 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10998__B net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09765_ net1098 game.CPU.applesa.ab.check_walls.above.walls\[97\] vssd1 vssd1 vccd1
+ vccd1 _04008_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout183_X net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Left_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11175__A game.CPU.applesa.ab.absxs.body_x\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_213_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09696_ net909 game.CPU.applesa.ab.absxs.body_y\[7\] game.CPU.applesa.ab.absxs.body_y\[5\]
+ net900 _03937_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__a221o_1
XANTENNA__17222__A1 _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_317_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14036__A1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14036__B2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1092_X net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_319_Left_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12047__B1 _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_239_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16981__B1 _02665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13795__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18594__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_340_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10540_ _03197_ _04606_ net754 vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__a21oi_4
XANTENNA__16194__D1 _02205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Left_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_269_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10471_ net929 net1268 vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12210_ game.CPU.applesa.ab.check_walls.above.walls\[173\] net548 vssd1 vssd1 vccd1
+ vccd1 _06096_ sky130_fd_sc_hd__xnor2_1
X_13190_ _07060_ _07061_ _07062_ _07063_ net498 net690 vssd1 vssd1 vccd1 vccd1 _07064_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_328_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12141_ net782 net552 vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_328_Left_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout96_X net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_285_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15764__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ game.CPU.applesa.ab.check_walls.above.walls\[85\] net386 vssd1 vssd1 vccd1
+ vccd1 _05959_ sky130_fd_sc_hd__nor2_1
Xhold590 game.writer.tracker.frame\[553\] vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_291_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11023_ game.CPU.applesa.ab.absxs.body_x\[91\] net546 vssd1 vssd1 vccd1 vccd1 _04913_
+ sky130_fd_sc_hd__xnor2_1
X_15900_ game.CPU.applesa.ab.absxs.body_y\[40\] net341 vssd1 vssd1 vccd1 vccd1 _01912_
+ sky130_fd_sc_hd__nand2_1
X_16880_ net135 _02272_ _02448_ _02632_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[258\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_218_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15831_ _03257_ net344 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_189_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14275__A1 game.CPU.applesa.ab.absxs.body_x\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19025__Q game.CPU.applesa.ab.check_walls.above.walls\[70\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ net602 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__inv_2
X_12974_ net508 _06847_ vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__or2_1
XFILLER_0_188_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15762_ game.CPU.applesa.ab.absxs.body_y\[117\] net446 vssd1 vssd1 vccd1 vccd1 _01774_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__13483__C1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_339_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17213__A1 _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17501_ _02778_ net427 _02841_ _02849_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__a31o_1
X_14713_ _03513_ _08547_ vssd1 vssd1 vccd1 vccd1 _08550_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_337_Left_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14027__A1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11925_ game.CPU.applesa.ab.check_walls.above.walls\[189\] net306 vssd1 vssd1 vccd1
+ vccd1 _05813_ sky130_fd_sc_hd__nor2_1
X_18481_ net636 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__inv_2
XFILLER_0_234_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18937__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15693_ _03248_ net350 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17432_ _02772_ _02825_ _02827_ _02861_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_123_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_346_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14644_ game.CPU.clock1.counter\[21\] _08484_ net268 vssd1 vssd1 vccd1 vccd1 _08485_
+ sky130_fd_sc_hd__o21ai_1
X_11856_ net804 net309 vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__nand2_1
XFILLER_0_345_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16972__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16882__Y _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10807_ game.CPU.applesa.ab.absxs.body_y\[18\] _04699_ _04700_ game.CPU.applesa.ab.absxs.body_y\[14\]
+ vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__a22o_1
X_14575_ game.CPU.clock1.counter\[20\] _03521_ game.CPU.speed1.Qa\[2\] vssd1 vssd1
+ vccd1 vccd1 _08437_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17363_ net1116 _02791_ _02792_ _02789_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__a22o_1
XANTENNA__15004__B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09454__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11787_ net574 _05254_ _05259_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09454__B2 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19102_ net1177 _00140_ _00773_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[147\]
+ sky130_fd_sc_hd__dfrtp_4
X_16314_ net1947 net720 _02304_ _02309_ _02273_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[14\]
+ sky130_fd_sc_hd__a32o_1
X_13526_ _07398_ _07399_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__and2_1
X_10738_ game.CPU.applesa.ab.absxs.body_y\[13\] _04653_ _04654_ game.CPU.applesa.ab.absxs.body_y\[9\]
+ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17294_ net2018 net722 _02755_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[549\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_55_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15939__B net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_250_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19033_ net1193 _00263_ _00704_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_13457_ net704 _07015_ _07330_ net512 vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__o211a_1
X_16245_ net244 _02227_ net222 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10669_ game.CPU.applesa.ab.absxs.body_x\[16\] _04699_ _04700_ game.CPU.applesa.ab.absxs.body_x\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__a22o_1
XANTENNA__13633__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12408_ game.CPU.applesa.ab.absxs.body_y\[54\] net521 net361 game.CPU.applesa.ab.absxs.body_y\[52\]
+ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15020__A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11013__B2 game.CPU.applesa.ab.absxs.body_x\[53\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_140_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13388_ _06870_ _06886_ net679 vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__mux2_1
X_16176_ _01854_ _01856_ _01859_ _01916_ _02187_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__o311a_1
XFILLER_0_267_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12339_ _04808_ _04220_ net1162 vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__mux2_1
X_15127_ net1208 net1233 game.CPU.applesa.ab.check_walls.above.walls\[155\] vssd1
+ vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__and3_1
XANTENNA__10164__A _03527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13893__A1_N net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18331__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_227_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19935_ clknet_leaf_38_clk game.writer.tracker.next_frame\[530\] net1325 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[530\] sky130_fd_sc_hd__dfrtp_1
X_15058_ net1211 net1237 net809 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__and3_1
XFILLER_0_282_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15674__B net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14009_ net876 game.CPU.applesa.ab.check_walls.above.walls\[139\] game.CPU.applesa.ab.check_walls.above.walls\[141\]
+ net861 _07881_ vssd1 vssd1 vccd1 vccd1 _07883_ sky130_fd_sc_hd__a221o_1
XFILLER_0_282_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_266_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19866_ clknet_leaf_20_clk game.writer.tracker.next_frame\[461\] net1310 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[461\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19712__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18817_ clknet_leaf_72_clk game.CPU.clock1.next_counter\[20\] _00554_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11707__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19797_ clknet_leaf_36_clk game.writer.tracker.next_frame\[392\] net1351 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[392\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_301_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09550_ net912 game.CPU.applesa.ab.absxs.body_x\[112\] game.CPU.applesa.ab.absxs.body_y\[114\]
+ net904 vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a22o_1
XANTENNA__15690__A game.CPU.applesa.ab.absxs.body_y\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18748_ clknet_leaf_64_clk _01165_ _00485_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_223_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17204__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09481_ net924 game.CPU.applesa.ab.check_walls.above.walls\[179\] _03478_ net1147
+ _03723_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__o221a_1
X_18679_ clknet_leaf_13_clk _01096_ _00416_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[117\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14018__A1 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_259_Right_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14018__B2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19862__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout143_A _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_195_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_351_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11252__B2 game.CPU.applesa.ab.absxs.body_x\[114\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15849__B net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_312_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout310_A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09847__B game.CPU.applesa.ab.absxs.body_y\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_332_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1052_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_310_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10763__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18241__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1317_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout311 net313 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__buf_4
XFILLER_0_273_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1309 net1314 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 net323 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_2
Xfanout333 game.CPU.walls.rand_wall.abduyd.next_wall\[6\] vssd1 vssd1 vccd1 vccd1
+ net333 sky130_fd_sc_hd__buf_4
Xfanout344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10515__B1 _04609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1105_X net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19392__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_323_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout366 net368 vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_4
XANTENNA__09381__B1 _03384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20006_ net1375 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XANTENNA__11617__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ net1083 _03278_ _03350_ net1146 vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__a22o_1
Xfanout377 net380 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_4
Xfanout388 net389 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_4
XANTENNA__14257__A1 game.CPU.applesa.ab.absxs.body_y\[76\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout944_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__buf_2
XANTENNA__14257__B2 game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_241_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09748_ _03985_ _03986_ _03989_ _03990_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout56_A _02354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10818__A1 game.CPU.applesa.ab.absxs.body_y\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09679_ net1111 game.CPU.applesa.ab.absxs.body_x\[100\] vssd1 vssd1 vccd1 vccd1 _03922_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__14009__A1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10818__B2 game.CPU.applesa.ab.absxs.body_y\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14009__B2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20011__A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09537__A1_N net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_226_Right_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11633__A game.CPU.applesa.ab.check_walls.above.walls\[157\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ _05379_ _05598_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.collision_leftn
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_87_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_328_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12690_ _06561_ _06563_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_327_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12448__B net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13768__B1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11641_ net564 _05525_ _05527_ _05529_ _05522_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10249__A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_343_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_Left_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_159_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16862__C _02608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14360_ net1266 net884 net873 net1265 vssd1 vssd1 vccd1 vccd1 _08234_ sky130_fd_sc_hd__o22a_1
X_11572_ game.CPU.applesa.ab.check_walls.above.walls\[129\] net769 vssd1 vssd1 vccd1
+ vccd1 _05461_ sky130_fd_sc_hd__xor2_1
XANTENNA__08942__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15759__B net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ net680 _06761_ _07184_ net204 vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__o211a_1
X_10523_ _04635_ game.CPU.applesa.ab.absxs.body_x\[61\] _04632_ vssd1 vssd1 vccd1
+ vccd1 _01180_ sky130_fd_sc_hd__mux2_1
XANTENNA__11794__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14291_ game.CPU.applesa.ab.absxs.body_x\[54\] net1056 vssd1 vssd1 vccd1 vccd1 _08165_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__12464__A game.CPU.applesa.ab.absxs.body_x\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09757__B game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13615__S0 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire756 _03526_ vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_122_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13242_ game.writer.tracker.frame\[504\] game.writer.tracker.frame\[505\] net1015
+ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__mux2_1
X_16030_ game.CPU.applesa.ab.absxs.body_x\[92\] net354 vssd1 vssd1 vccd1 vccd1 _02042_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_220_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10454_ net850 _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__nor2_2
XFILLER_0_296_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13173_ _06984_ _07046_ net177 vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__a21o_1
X_10385_ net1125 game.CPU.apple_location\[7\] vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_248_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12124_ game.CPU.applesa.ab.check_walls.above.walls\[175\] net295 net289 game.CPU.applesa.ab.check_walls.above.walls\[174\]
+ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__o22a_1
XANTENNA__16485__A2 _02432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19735__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_248_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_264_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17981_ net606 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_53_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_261_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_155_Left_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19720_ clknet_leaf_35_clk game.writer.tracker.next_frame\[315\] net1346 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[315\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_248_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_236_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16932_ _02364_ net87 _02651_ net1596 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[291\]
+ sky130_fd_sc_hd__a22o_1
X_12055_ _05939_ _05940_ _05941_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__or3_1
XFILLER_0_263_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16237__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ _03307_ net543 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_183_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17434__A1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19651_ clknet_leaf_21_clk game.writer.tracker.next_frame\[246\] net1342 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[246\] sky130_fd_sc_hd__dfrtp_1
X_16863_ net1473 _02626_ _02627_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[246\]
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_125_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14248__B2 game.CPU.applesa.ab.absxs.body_y\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16788__A3 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19885__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18602_ clknet_leaf_65_clk _01022_ _00339_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[83\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_345_Left_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15814_ _01815_ _01816_ _01819_ _01822_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__or4_1
X_19582_ clknet_leaf_34_clk game.writer.tracker.next_frame\[177\] net1349 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[177\] sky130_fd_sc_hd__dfrtp_1
X_16794_ _02472_ net102 _02599_ net1584 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[205\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18533_ net629 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__inv_2
XANTENNA__10809__A1 game.CPU.applesa.ab.absxs.body_y\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_232_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15745_ _03469_ net269 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10809__B2 game.CPU.applesa.ab.absxs.body_y\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12957_ net505 _06830_ _06829_ net205 vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11543__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15015__A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18464_ net652 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__inv_2
XANTENNA__11482__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11908_ net750 _05283_ _05795_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_259_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ _03383_ net473 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__nand2_1
X_12888_ game.writer.tracker.frame\[64\] game.writer.tracker.frame\[65\] net1039 vssd1
+ vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__mux2_2
XFILLER_0_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_358_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12358__B net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_164_Left_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_272_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13759__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17415_ _02779_ _02842_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__nor2_1
XANTENNA__09013__A game.CPU.applesa.ab.absxs.body_x\[96\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14627_ _08474_ net267 _08473_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[14\]
+ sky130_fd_sc_hd__and3b_1
X_11839_ net747 _05429_ _05431_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__o21ai_1
X_18395_ net619 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18326__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14420__B2 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17346_ _02773_ _02775_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14558_ net453 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.abduyd.next_wall\[4\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__15669__B net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12431__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_333_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12982__A1 _06852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19265__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_354_Left_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13509_ net511 _07301_ _07303_ net228 vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17277_ _02259_ _02421_ _02750_ net1994 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[537\]
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13606__S0 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14489_ _08078_ _08081_ _08062_ vssd1 vssd1 vccd1 vccd1 _08363_ sky130_fd_sc_hd__o21a_1
XANTENNA__16712__A3 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19016_ net1195 _00245_ _00687_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[61\]
+ sky130_fd_sc_hd__dfrtp_4
X_16228_ net177 net141 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__or2_4
XFILLER_0_3_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_341_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12093__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12734__A1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12661__X _06538_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16159_ _01711_ _01712_ _01903_ _02151_ _02170_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_173_Left_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08981_ game.CPU.applesa.ab.absxs.body_x\[93\] vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_283_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_328_Right_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13409__S net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_225_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19918_ clknet_leaf_33_clk game.writer.tracker.next_frame\[513\] net1301 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[513\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_299_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17425__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19849_ clknet_leaf_37_clk game.writer.tracker.next_frame\[444\] net1356 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[444\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09902__A2 _03684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09602_ net1101 game.CPU.applesa.ab.absxs.body_x\[73\] vssd1 vssd1 vccd1 vccd1 _03845_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_155_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09533_ net1098 game.CPU.applesa.ab.check_walls.above.walls\[73\] vssd1 vssd1 vccd1
+ vccd1 _03776_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout260_A net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_182_Left_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_305_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ net906 net1172 _03705_ _03706_ net1263 vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_309_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12268__B net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19608__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_236_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09395_ _03635_ _03636_ _03637_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__or3_4
XANTENNA__12836__X _06710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout525_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14411__A1 game.CPU.applesa.ab.absxs.body_x\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout146_X net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18236__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16149__D1 _01618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__B1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15579__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10579__A3 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1055_X net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14175__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18632__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19758__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13073__S1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout894_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_191_Left_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13667__X _07541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13922__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_325_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09593__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10170_ net1134 _04362_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_301_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16978__X _02665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14478__A1 game.CPU.applesa.ab.absxs.body_y\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_266_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14478__B2 game.CPU.applesa.ab.absxs.body_y\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18782__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1106 net1108 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_8
Xfanout1117 game.CPU.bodymain1.main.score\[3\] vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__clkbuf_2
Xfanout130 _02276_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10532__A _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_245_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_6_0_clk_X clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1128 net1129 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__clkbuf_8
Xfanout141 _02231_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15734__A2_N net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1139 net1143 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__buf_6
Xfanout152 net155 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09880__X _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_233_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout163 net164 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__buf_2
Xfanout174 _06702_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout185 net187 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10251__B _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout947_X net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 _02289_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_4
X_13860_ game.writer.tracker.frame\[555\] net708 net671 game.writer.tracker.frame\[556\]
+ _07733_ vssd1 vssd1 vccd1 vccd1 _07734_ sky130_fd_sc_hd__o221a_1
XFILLER_0_214_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19138__CLK net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout59_X net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12811_ game.writer.tracker.frame\[366\] game.writer.tracker.frame\[367\] net997
+ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__mux2_1
XANTENNA__13989__B1 game.CPU.applesa.ab.check_walls.above.walls\[21\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13791_ game.writer.tracker.frame\[425\] game.writer.tracker.frame\[427\] game.writer.tracker.frame\[428\]
+ game.writer.tracker.frame\[426\] net977 net1020 vssd1 vssd1 vccd1 vccd1 _07665_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_336_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13054__S net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15530_ net888 net1057 _01551_ _01508_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__a31o_1
XFILLER_0_198_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12742_ game.writer.tracker.frame\[66\] game.writer.tracker.frame\[67\] net1026 vssd1
+ vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__mux2_1
XANTENNA__16927__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19288__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12893__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20051__1369 vssd1 vssd1 vccd1 vccd1 _20051__1369/HI net1369 sky130_fd_sc_hd__conb_1
X_12673_ _03363_ game.writer.updater.commands.mode\[1\] game.writer.updater.commands.mode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__or3b_1
X_15461_ _01450_ _01462_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12746__X _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__Y _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_315_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17200_ _02509_ net71 net716 vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__o21a_1
XANTENNA__12379__A1_N game.CPU.applesa.ab.absxs.body_y\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_182_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11624_ _05512_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__inv_2
X_14412_ game.CPU.applesa.ab.absxs.body_x\[46\] net878 net864 game.CPU.applesa.ab.absxs.body_y\[45\]
+ vssd1 vssd1 vccd1 vccd1 _08286_ sky130_fd_sc_hd__a2bb2o_1
X_18180_ net608 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__inv_2
XANTENNA__09768__A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15392_ _03363_ _03364_ game.writer.updater.commands.mode\[0\] vssd1 vssd1 vccd1
+ vccd1 _08934_ sky130_fd_sc_hd__and3_2
XFILLER_0_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_331_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12964__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17131_ _02390_ net76 _02712_ net1917 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[429\]
+ sky130_fd_sc_hd__a22o_1
X_11555_ game.CPU.applesa.ab.check_walls.above.walls\[192\] net775 vssd1 vssd1 vccd1
+ vccd1 _05444_ sky130_fd_sc_hd__xor2_1
X_14343_ _03245_ net1063 net878 game.CPU.applesa.ab.absxs.body_x\[38\] _08214_ vssd1
+ vssd1 vccd1 vccd1 _08217_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ _04156_ _04607_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__nand2_8
XFILLER_0_135_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17062_ net189 net173 _02229_ net717 vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__o31a_2
X_14274_ game.CPU.applesa.ab.absxs.body_x\[49\] net883 net874 game.CPU.applesa.ab.absxs.body_x\[51\]
+ _08147_ vssd1 vssd1 vccd1 vccd1 _08148_ sky130_fd_sc_hd__o221a_1
XFILLER_0_122_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11486_ net819 net256 _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15001__C game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_311_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11519__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13225_ _07096_ _07097_ net690 vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__mux2_1
X_16013_ _03239_ net351 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13913__B1 game.CPU.applesa.ab.check_walls.above.walls\[124\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10437_ game.CPU.applesa.ab.absxs.body_x\[4\] _04156_ net754 net1438 vssd1 vssd1
+ vccd1 vccd1 _01207_ sky130_fd_sc_hd__o22a_1
XANTENNA__17104__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_296_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13156_ net705 _07029_ _07026_ net231 vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_131_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ game.CPU.applesa.ab.absxs.body_y\[5\] net848 _04158_ net1445 vssd1 vssd1
+ vccd1 vccd1 _01274_ sky130_fd_sc_hd__a22o_1
XFILLER_0_237_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16113__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12107_ net818 net296 vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__nand2_1
X_13087_ game.writer.tracker.frame\[202\] game.writer.tracker.frame\[203\] net1011
+ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__mux2_1
X_17964_ net658 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__inv_2
X_10299_ net1264 game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__nand2b_4
X_19703_ clknet_leaf_30_clk game.writer.tracker.next_frame\[298\] net1284 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[298\] sky130_fd_sc_hd__dfrtp_1
X_16915_ _02335_ _02644_ net728 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__o21a_1
X_12038_ game.CPU.applesa.ab.check_walls.above.walls\[143\] net293 net288 net791 vssd1
+ vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__15952__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17895_ net643 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__inv_2
XANTENNA__13692__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11152__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19634_ clknet_leaf_28_clk game.writer.tracker.next_frame\[229\] net1290 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[229\] sky130_fd_sc_hd__dfrtp_1
X_16846_ _02520_ net98 _02619_ net717 vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__o31a_1
XANTENNA__13429__C1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16630__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19565_ clknet_leaf_34_clk game.writer.tracker.next_frame\[160\] net1333 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[160\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_220_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16777_ _02443_ net109 _02594_ game.writer.tracker.frame\[193\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[193\] sky130_fd_sc_hd__a22o_1
XANTENNA__19213__Q game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13989_ net884 game.CPU.applesa.ab.check_walls.above.walls\[17\] game.CPU.applesa.ab.check_walls.above.walls\[21\]
+ net864 _07859_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_245_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18516_ net583 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__inv_2
X_15728_ game.CPU.applesa.ab.absxs.body_x\[12\] net355 vssd1 vssd1 vccd1 vccd1 _01740_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19496_ clknet_leaf_25_clk game.writer.tracker.next_frame\[91\] net1321 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[91\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_272_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12652__B1 game.CPU.applesa.twoapples.absxs.next_head\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_18447_ net592 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15659_ game.CPU.applesa.ab.check_walls.above.walls\[48\] net273 vssd1 vssd1 vccd1
+ vccd1 _01671_ sky130_fd_sc_hd__or2_1
XFILLER_0_307_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18655__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09180_ net806 vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__inv_2
X_18378_ net600 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_192_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19900__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17329_ _02275_ _02435_ _02764_ net1850 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[575\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_231_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload45_A clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13928__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__B1 _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout106_A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_287_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13380__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_255_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12551__B net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17110__A3 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13139__S net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16023__B net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11448__A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ game.CPU.applesa.ab.start_enable vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__inv_2
XFILLER_0_227_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15862__B net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_320_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_270_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_316_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09639__A1 net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19430__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12279__A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09639__B2 net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09516_ net1159 game.CPU.applesa.ab.absxs.body_y\[48\] vssd1 vssd1 vccd1 vccd1 _03759_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__11446__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09447_ net920 game.CPU.applesa.ab.check_walls.above.walls\[138\] game.CPU.applesa.ab.check_walls.above.walls\[141\]
+ net897 vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_26_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_332_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14494__A _08362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13818__S0 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout907_A _03199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13199__A1 game.writer.tracker.frame\[401\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09378_ net916 game.CPU.applesa.ab.check_walls.above.walls\[9\] game.CPU.applesa.ab.check_walls.above.walls\[12\]
+ net893 _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19580__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12946__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12726__B net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_331_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09875__X _04118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11340_ net743 _05226_ _05228_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_132_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16688__A2 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_269_Left_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ _04831_ _05031_ _05152_ _05160_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__and4_1
XFILLER_0_132_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16214__A _02163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13010_ game.writer.tracker.frame\[516\] game.writer.tracker.frame\[517\] net1008
+ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__mux2_1
X_10222_ _04404_ _04414_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__or2_1
XANTENNA__12174__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12461__B net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_246_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_245_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15648__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11358__A game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _04347_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__inv_2
XANTENNA__16860__A2 _02412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14320__B1 net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11077__B net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15772__B net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ _04290_ _04291_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__xnor2_1
X_14961_ _08699_ _08737_ _08659_ vssd1 vssd1 vccd1 vccd1 _08738_ sky130_fd_sc_hd__a21o_1
Xhold8 game.CPU.left_button.sync1.Q vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ net63 _02566_ net559 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_233_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13912_ net867 game.CPU.applesa.ab.check_walls.above.walls\[124\] game.CPU.applesa.ab.check_walls.above.walls\[122\]
+ net877 vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12882__A0 _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17680_ game.CPU.walls.rand_wall.count_luck\[2\] game.CPU.walls.rand_wall.count_luck\[1\]
+ _03063_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__and3_1
XANTENNA__14021__X _07895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10488__A2 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14892_ _08659_ _08662_ _08665_ _08668_ vssd1 vssd1 vccd1 vccd1 _08669_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_278_Left_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16631_ _02237_ _02302_ _02517_ net713 vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__o31a_1
X_13843_ game.writer.tracker.frame\[526\] net842 net708 game.writer.tracker.frame\[527\]
+ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__o22a_1
XANTENNA__12189__A net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15820__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19350_ clknet_leaf_70_clk game.CPU.applesa.twoapples.absxs.next_head\[6\] vssd1
+ vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.y_final\[2\] sky130_fd_sc_hd__dfxtp_1
XANTENNA__11437__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16562_ net154 _02327_ net127 _02488_ net1666 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[84\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__18678__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13774_ game.writer.tracker.frame\[153\] net838 net674 game.writer.tracker.frame\[156\]
+ vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__o22a_1
X_10986_ _03322_ net401 vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19923__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18301_ net641 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_256_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15513_ _01518_ _01530_ _01535_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__and3_1
XFILLER_0_328_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12725_ net841 net840 vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__and2_1
X_19281_ clknet_leaf_67_clk _01330_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.count\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16493_ net183 net167 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__nor2_2
XFILLER_0_242_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13809__S0 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18232_ net665 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
X_15444_ _08903_ _08922_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_178_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_242_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12656_ game.CPU.applesa.ab.absxs.body_x\[66\] net373 net530 game.CPU.applesa.ab.absxs.body_x\[67\]
+ _06532_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__o221a_1
XANTENNA__10660__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18163_ net583 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__inv_2
XANTENNA__11540__B net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11607_ net568 _05489_ _05493_ _05494_ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__a2111o_1
XANTENNA__15012__B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17325__B1 _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15375_ _08885_ _08916_ vssd1 vssd1 vccd1 vccd1 _08917_ sky130_fd_sc_hd__nand2_1
XANTENNA__16128__B2 game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12587_ game.CPU.applesa.ab.absxs.body_y\[89\] net523 vssd1 vssd1 vccd1 vccd1 _06464_
+ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_287_Left_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17114_ net158 net66 net80 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__and3_1
X_14326_ game.CPU.applesa.ab.absxs.body_y\[75\] net941 vssd1 vssd1 vccd1 vccd1 _08200_
+ sky130_fd_sc_hd__nand2_1
X_11538_ game.CPU.applesa.ab.check_walls.above.walls\[144\] net773 vssd1 vssd1 vccd1
+ vccd1 _05427_ sky130_fd_sc_hd__xnor2_1
X_18094_ net606 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15947__B net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold408 game.writer.tracker.frame\[40\] vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold419 game.writer.tracker.frame\[344\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
X_17045_ _02542_ net88 _02684_ net1614 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[371\]
+ sky130_fd_sc_hd__a22o_1
X_14257_ game.CPU.applesa.ab.absxs.body_y\[76\] net869 net854 game.CPU.applesa.ab.absxs.body_y\[78\]
+ _08130_ vssd1 vssd1 vccd1 vccd1 _08131_ sky130_fd_sc_hd__a221o_1
X_11469_ game.CPU.applesa.ab.check_walls.above.walls\[21\] net318 _05356_ _05357_
+ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19303__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ game.writer.tracker.frame\[430\] game.writer.tracker.frame\[431\] net1020
+ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_267_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14188_ _08055_ _08057_ _08059_ _08061_ vssd1 vssd1 vccd1 vccd1 _08062_ sky130_fd_sc_hd__or4_2
XANTENNA__12371__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19208__Q game.CPU.applesa.ab.YMAX\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_280_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ _07007_ _07012_ net224 vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10172__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18996_ net1194 _00223_ _00667_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[41\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_264_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13114__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09961__A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15682__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17947_ net639 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__inv_2
XANTENNA__09869__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_296_Left_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19453__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09869__B2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11676__A1 game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09680__B game.CPU.applesa.ab.absxs.body_x\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17878_ net656 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__inv_2
XFILLER_0_252_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16603__A2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17800__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19617_ clknet_leaf_21_clk game.writer.tracker.next_frame\[212\] net1336 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[212\] sky130_fd_sc_hd__dfrtp_1
X_16829_ net1741 _02610_ _02611_ net132 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[228\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_356_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12099__A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19548_ clknet_leaf_49_clk game.writer.tracker.next_frame\[143\] net1279 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[143\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10111__S _04311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_278_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09301_ _03533_ _03534_ _03540_ _03541_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18782__Q game.CPU.applesa.ab.absxs.body_x\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13930__B net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19479_ clknet_leaf_18_clk game.writer.tracker.next_frame\[74\] net1315 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[74\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17402__B game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12827__A net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17564__B1 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09232_ net782 vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__inv_2
XANTENNA__14378__B1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_233_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12928__A1 _06795_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16018__B net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12928__B2 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16119__A1 game.CPU.applesa.ab.check_walls.above.walls\[177\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ game.CPU.applesa.ab.check_walls.above.walls\[58\] vssd1 vssd1 vccd1 vccd1
+ _03412_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout223_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16119__B2 game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15590__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18514__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09094_ game.CPU.applesa.ab.absxs.body_y\[42\] vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09855__B game.CPU.applesa.ab.absxs.body_y\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout109_X net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_309_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16034__A game.CPU.applesa.ab.absxs.body_x\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1132_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_247_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15873__A game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11903__A2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17095__A2 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09996_ net2031 net1996 _04207_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__mux2_1
XANTENNA__09871__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18957__Q game.CPU.applesa.ab.check_walls.above.walls\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08947_ net1117 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Left_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12313__C1 _06198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout857_A _03376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11906__A game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_270_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19946__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11625__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13680__X _07554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_300_Left_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11419__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10840_ _03511_ game.CPU.randy.counter1.count\[4\] game.CPU.randy.counter1.count\[3\]
+ _03513_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_333_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18692__Q game.CPU.applesa.ab.absxs.body_x\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12040__A2_N net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ game.CPU.applesa.ab.absxs.body_y\[73\] _04675_ _04676_ game.CPU.applesa.ab.absxs.body_y\[69\]
+ vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__a22o_1
X_12510_ game.CPU.applesa.ab.absxs.body_x\[72\] net384 vssd1 vssd1 vccd1 vccd1 _06387_
+ sky130_fd_sc_hd__xnor2_1
X_13490_ net508 _07123_ net700 vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__a21o_1
XFILLER_0_353_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12441_ game.CPU.applesa.ab.absxs.body_x\[105\] net378 net361 game.CPU.applesa.ab.absxs.body_y\[104\]
+ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__o22a_1
XFILLER_0_191_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_22_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10257__A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19326__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12395__A2 game.CPU.applesa.twoapples.absxs.next_head\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12372_ game.CPU.applesa.ab.absxs.body_x\[114\] net372 vssd1 vssd1 vccd1 vccd1 _06249_
+ sky130_fd_sc_hd__xnor2_1
X_15160_ net1213 net1239 net782 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__and3_1
XFILLER_0_288_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_251_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08950__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14111_ net947 game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1 vccd1
+ vccd1 _07985_ sky130_fd_sc_hd__xor2_1
X_11323_ net563 _04775_ game.CPU.applesa.ab.apple_possible\[5\] vssd1 vssd1 vccd1
+ vccd1 _05212_ sky130_fd_sc_hd__o21ai_1
X_15091_ net1211 net1237 net796 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__and3_1
XFILLER_0_278_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_37_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14042_ net885 net874 _06549_ vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__and3_1
X_11254_ game.CPU.applesa.ab.absxs.body_x\[111\] net545 net539 game.CPU.applesa.ab.absxs.body_y\[110\]
+ _05132_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__a221o_1
XANTENNA__19476__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19028__Q game.CPU.applesa.ab.check_walls.above.walls\[73\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _04386_ _04387_ _04385_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__a21o_1
XANTENNA__17086__A2 _02479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18850_ clknet_leaf_6_clk _01241_ _00560_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_11185_ game.CPU.applesa.ab.absxs.body_y\[86\] net403 vssd1 vssd1 vccd1 vccd1 _05075_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17801_ _03138_ _03139_ net992 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__mux2_1
XANTENNA__16833__A2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10136_ game.CPU.randy.f1.c1.count\[6\] game.CPU.randy.f1.c1.count\[9\] game.CPU.randy.f1.c1.count\[8\]
+ game.CPU.randy.f1.c1.count\[11\] vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__or4_1
X_18781_ clknet_leaf_63_clk _01198_ _00518_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[95\]
+ sky130_fd_sc_hd__dfrtp_4
X_15993_ game.CPU.applesa.ab.check_walls.above.walls\[98\] net469 vssd1 vssd1 vccd1
+ vccd1 _02005_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14399__A game.CPU.applesa.ab.absxs.body_y\[69\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_206_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17732_ net1912 _03097_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__xnor2_1
X_10067_ _04223_ _04274_ _04238_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__a21o_1
X_14944_ _08711_ _08720_ vssd1 vssd1 vccd1 vccd1 _08721_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11658__A1 game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11658__B2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17663_ net1753 _03052_ _03054_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11535__B net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15007__B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14875_ game.CPU.walls.abc.number\[7\] game.CPU.walls.abc.number\[3\] game.CPU.walls.abc.counter
+ vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__mux2_1
X_19402_ clknet_leaf_47_clk _01402_ net1279 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.x\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkload1_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16614_ net206 _02266_ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__nor2_4
XANTENNA__17062__X _02689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13826_ _07620_ _07699_ net174 vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__a21o_1
X_17594_ _03009_ _03012_ net582 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19333_ clknet_leaf_71_clk _01349_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.count_luck\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_16545_ net1714 _02474_ _02476_ net124 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[79\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13757_ game.writer.tracker.frame\[135\] net708 net671 game.writer.tracker.frame\[136\]
+ vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__o22a_1
X_10969_ game.CPU.applesa.ab.absxs.body_y\[101\] net404 vssd1 vssd1 vccd1 vccd1 _04859_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__17010__A2 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12708_ _06565_ _06581_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__nor2_1
XANTENNA__10633__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19264_ clknet_leaf_8_clk _00052_ _00894_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11291__C1 _04894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16476_ _02289_ _02385_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__nand2_4
XFILLER_0_72_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13688_ _07558_ _07561_ net221 vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18215_ net666 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__inv_2
XFILLER_0_316_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15427_ _01449_ _01454_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19195_ clknet_leaf_54_clk net334 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.y_final\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12639_ game.CPU.applesa.ab.absxs.body_x\[19\] net531 net519 game.CPU.applesa.ab.absxs.body_y\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__a22o_1
XANTENNA__18334__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18146_ net626 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__inv_2
XFILLER_0_331_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15358_ _08885_ _08898_ vssd1 vssd1 vccd1 vccd1 _08900_ sky130_fd_sc_hd__or2_1
XFILLER_0_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15677__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_269_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_215_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13478__A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire180 net181 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_2
Xhold205 game.writer.tracker.frame\[299\] vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
X_14309_ _08179_ _08180_ _08175_ _08177_ vssd1 vssd1 vccd1 vccd1 _08183_ sky130_fd_sc_hd__a211o_1
XANTENNA__19819__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_300_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18077_ net669 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__inv_2
XANTENNA__09675__B net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold216 game.writer.tracker.frame\[430\] vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ _08815_ _08837_ _08839_ _08817_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a22o_1
Xhold227 game.writer.tracker.frame\[496\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 game.writer.tracker.frame\[443\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_wire181_X net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold249 game.writer.tracker.frame\[86\] vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ _02369_ net85 _02680_ net1625 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[358\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17077__A2 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout707 _06599_ vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_4
X_09850_ net1134 game.CPU.applesa.ab.absxs.body_y\[30\] vssd1 vssd1 vccd1 vccd1 _04093_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_70_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout718 net719 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_113_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 net731 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_265_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09691__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09781_ net1089 _03457_ net790 net892 _04020_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__a221o_1
X_18979_ net1201 _00204_ _00650_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_304_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19587__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14102__A net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_240_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout173_A _06702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18509__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13941__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12828__Y _06702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19401__Q game.CPU.applesa.x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1082_A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_313_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout438_A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19349__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10624__A2 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_315_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09215_ game.CPU.applesa.ab.check_walls.above.walls\[160\] vssd1 vssd1 vccd1 vccd1
+ _03464_ sky130_fd_sc_hd__inv_2
XANTENNA__11180__B net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16760__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10077__A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout226_X net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout605_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1347_A net1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09866__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12377__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ net825 vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__inv_2
XFILLER_0_350_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10388__A1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15587__B net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19499__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09077_ game.CPU.applesa.ab.absxs.body_y\[90\] vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__inv_2
XANTENNA__16512__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12292__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1135_X net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_303_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14523__B1 _07164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_275_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout974_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_338_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1302_X net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11888__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11888__B2 game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout86_A _02638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_338_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16815__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_256_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ _04204_ _04205_ _04159_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_274_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12990_ game.writer.tracker.frame\[550\] game.writer.tracker.frame\[551\] net1006
+ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__mux2_1
XANTENNA__14012__A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16028__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_271_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11355__B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11941_ _05822_ _05823_ _05827_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__and4_1
XANTENNA__16579__A1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17240__A2 _02432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14660_ _08490_ net266 vssd1 vssd1 vccd1 vccd1 _08499_ sky130_fd_sc_hd__or2_1
X_11872_ net831 net312 _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08945__A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13611_ game.writer.tracker.frame\[261\] game.writer.tracker.frame\[263\] game.writer.tracker.frame\[264\]
+ game.writer.tracker.frame\[262\] net967 net996 vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__mux4_1
XANTENNA__12065__A1 game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10823_ _04482_ _04563_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__nor2_1
X_14591_ game.CPU.clock1.counter\[0\] net268 vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[0\]
+ sky130_fd_sc_hd__and2b_1
XANTENNA__12065__B2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12467__A game.CPU.applesa.ab.absxs.body_x\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13801__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_223_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11371__A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16330_ _02274_ _02322_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_253_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13542_ _07414_ _07415_ net488 vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11812__A1 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10615__A2 _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10754_ game.CPU.applesa.ab.absxs.body_y\[109\] _04665_ _04666_ game.CPU.applesa.ab.absxs.body_y\[105\]
+ vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11812__B2 game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12186__B net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09481__A2 game.CPU.applesa.ab.check_walls.above.walls\[179\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_299_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16881__B net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16200__B1 net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11090__B net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ net225 _02266_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__nor2_8
XANTENNA__15778__A game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_175_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18716__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13473_ _07076_ _07096_ net684 vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__mux2_1
X_10685_ _04593_ net329 vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16226__X _02234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_353_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18000_ net637 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__inv_2
X_15212_ game.CPU.applesa.normal1.number\[3\] _08773_ vssd1 vssd1 vccd1 vccd1 _08779_
+ sky130_fd_sc_hd__nand2_1
X_12424_ _06293_ _06295_ _06299_ _06300_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__or4b_1
X_16192_ _01879_ _01880_ _02200_ _02203_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_341_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10379__A1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15143_ net1210 net1236 game.CPU.applesa.ab.check_walls.above.walls\[171\] vssd1
+ vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__and3_1
X_12355_ _03236_ game.CPU.applesa.twoapples.absxs.next_head\[1\] vssd1 vssd1 vccd1
+ vccd1 _06232_ sky130_fd_sc_hd__nor2_1
XANTENNA__09495__B net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13317__A1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14514__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ game.CPU.applesa.ab.apple_possible\[7\] _05194_ vssd1 vssd1 vccd1 vccd1 _05195_
+ sky130_fd_sc_hd__xnor2_2
XFILLER_0_294_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19951_ clknet_leaf_43_clk game.writer.tracker.next_frame\[546\] net1307 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[546\] sky130_fd_sc_hd__dfrtp_1
X_12286_ game.CPU.applesa.ab.check_walls.above.walls\[135\] net422 vssd1 vssd1 vccd1
+ vccd1 _06172_ sky130_fd_sc_hd__nor2_1
X_15074_ net1216 net1238 net803 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__and3_1
XFILLER_0_278_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_264_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_248_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11237_ _05119_ _05120_ _05121_ _05126_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__or4_1
X_14025_ net984 game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1 vccd1
+ vccd1 _07899_ sky130_fd_sc_hd__xor2_1
X_18902_ clknet_leaf_4_clk _01269_ _00586_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11879__A1 game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19882_ clknet_leaf_26_clk game.writer.tracker.next_frame\[477\] net1319 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[477\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11879__B2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16402__A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16806__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_248_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18597__Q game.CPU.applesa.ab.absxs.body_y\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_18833_ clknet_leaf_0_clk _01224_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_11168_ game.CPU.applesa.ab.absxs.body_y\[76\] net534 vssd1 vssd1 vccd1 vccd1 _05058_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_186_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11546__A game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ _04319_ net1448 _04311_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18764_ clknet_leaf_51_clk _01181_ _00501_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[62\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15018__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11099_ game.CPU.applesa.ab.absxs.body_y\[56\] net536 vssd1 vssd1 vccd1 vccd1 _04989_
+ sky130_fd_sc_hd__nand2_1
X_15976_ _01981_ _01982_ _01983_ _01986_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__or4_1
X_17715_ net1574 _03084_ _03087_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__o21a_1
XANTENNA__15960__B game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14927_ _08662_ _08702_ vssd1 vssd1 vccd1 vccd1 _08704_ sky130_fd_sc_hd__xnor2_1
X_18695_ clknet_leaf_59_clk _01112_ _00432_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[41\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__18329__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13761__A net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17646_ game.CPU.kyle.L1.cnt_500hz\[6\] _08804_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_353_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14858_ net1816 _08647_ vssd1 vssd1 vccd1 vccd1 _08650_ sky130_fd_sc_hd__nor2_1
XFILLER_0_348_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12577__A2_N net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13809_ game.writer.tracker.frame\[441\] game.writer.tracker.frame\[443\] game.writer.tracker.frame\[444\]
+ game.writer.tracker.frame\[442\] net980 net1040 vssd1 vssd1 vccd1 vccd1 _07683_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17577_ net1440 net264 _02871_ _08809_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_275_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14789_ game.CPU.randy.counter1.count\[4\] _08604_ net138 vssd1 vssd1 vccd1 vccd1
+ _08607_ sky130_fd_sc_hd__o21ai_1
X_19316_ clknet_leaf_71_clk _01340_ _00922_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.apple_location2_n\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_325_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16528_ _02298_ _02376_ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__nor2_4
XFILLER_0_329_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_217_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_280_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19247_ clknet_leaf_17_clk _00061_ _00885_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15688__A game.CPU.applesa.ab.absxs.body_y\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16459_ net117 net166 _02415_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_139_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_304_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19641__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16742__A1 _02382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16136__X _02148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_317_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18064__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09000_ game.CPU.applesa.ab.absxs.body_x\[22\] vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__inv_2
Xclkbuf_3_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_332_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19178_ clknet_leaf_6_clk _01297_ _00840_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_289_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18129_ net578 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__inv_2
XFILLER_0_332_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_289_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13308__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14505__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19791__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10790__A1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_286_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13859__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09902_ _03677_ _03684_ _04143_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__o211a_1
XFILLER_0_300_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17408__A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout504 net516 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_228_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout515 net516 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_300_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12531__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20022_ net1276 vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
Xfanout526 net527 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_4
X_09833_ net923 game.CPU.applesa.ab.absxs.body_x\[106\] game.CPU.applesa.ab.absxs.body_x\[104\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__o22a_1
Xfanout537 game.CPU.applesa.ab.absxs.next_head\[4\] vssd1 vssd1 vccd1 vccd1 net537
+ sky130_fd_sc_hd__buf_4
Xfanout548 net550 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_4
Xfanout559 net560 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__buf_4
XANTENNA_fanout290_A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_207_Right_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16031__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__B2 game.CPU.applesa.ab.absxs.body_x\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ net898 net804 vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_308_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_253_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11175__B net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15870__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09695_ net1130 _03215_ _03216_ net1148 _03936_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout176_X net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18239__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1297_A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17222__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19171__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_317_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14036__A2 game.CPU.applesa.ab.check_walls.above.walls\[113\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16430__B1 _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_355_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18739__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16981__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout722_A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19131__Q game.CPU.applesa.ab.check_walls.above.walls\[176\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_239_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1085_X net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16733__A1 _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18889__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09596__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10470_ _04592_ _04600_ _04589_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_340_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_269_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09129_ game.CPU.applesa.ab.check_walls.above.walls\[0\] vssd1 vssd1 vccd1 vccd1
+ _03378_ sky130_fd_sc_hd__inv_2
XANTENNA__14007__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16497__B1 _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_328_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12140_ _05507_ _05508_ _05510_ _05512_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__or4_1
XFILLER_0_349_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_276_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout977_X net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ game.CPU.applesa.ab.check_walls.above.walls\[85\] _05192_ _05863_ vssd1 vssd1
+ vccd1 vccd1 _05958_ sky130_fd_sc_hd__and3_1
XANTENNA__17318__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold580 game.writer.tracker.frame\[16\] vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_285_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold591 game.CPU.walls.rand_wall.count_luck\[5\] vssd1 vssd1 vccd1 vccd1 net1976
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout89_X net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11022_ _03327_ net533 vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_263_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11366__A game.CPU.applesa.ab.check_walls.above.walls\[34\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15830_ _03284_ net355 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__nand2_1
XFILLER_0_218_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19514__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14275__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11085__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15761_ _03287_ net351 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_51_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ _06641_ _06643_ net686 vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__mux2_1
XANTENNA__12896__S net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17500_ _02825_ net426 _02840_ _02928_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_339_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17213__A2 net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10420__D _04563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14712_ _08548_ vssd1 vssd1 vccd1 vccd1 _08549_ sky130_fd_sc_hd__inv_2
X_11924_ net782 net391 net300 game.CPU.applesa.ab.check_walls.above.walls\[190\] vssd1
+ vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__o22a_1
X_18480_ net635 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__inv_2
X_15692_ game.CPU.applesa.ab.absxs.body_x\[28\] net354 vssd1 vssd1 vccd1 vccd1 _01704_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_231_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14396__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17431_ net1275 game.CPU.speed1.Qa\[0\] _02782_ net427 vssd1 vssd1 vccd1 vccd1 _02861_
+ sky130_fd_sc_hd__o211a_1
X_14643_ _08484_ net268 _08483_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[20\]
+ sky130_fd_sc_hd__and3b_1
XANTENNA__17988__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12038__B2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11855_ net804 net309 vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__or2_1
XANTENNA__19664__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15775__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12197__A net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_345_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13786__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12589__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13330__S0 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17362_ _02789_ _02790_ _02791_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__a21oi_2
X_10806_ game.CPU.applesa.ab.absxs.body_y\[19\] _04699_ _04700_ game.CPU.applesa.ab.absxs.body_y\[15\]
+ vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__a22o_1
X_14574_ net1275 _03519_ _08435_ game.CPU.clock1.counter\[1\] game.CPU.clock1.counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08436_ sky130_fd_sc_hd__a2111o_1
XANTENNA__15004__C game.CPU.applesa.ab.check_walls.above.walls\[32\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11786_ net823 net309 vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__xnor2_1
X_19101_ net1177 _00139_ _00772_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[146\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16313_ net196 _02308_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__nor2_4
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13525_ _06703_ _07253_ _07257_ _07289_ net162 vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__o32a_2
X_17293_ net130 _02365_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__or2_1
XFILLER_0_250_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10737_ game.CPU.applesa.ab.absxs.body_y\[14\] _04653_ _04654_ game.CPU.applesa.ab.absxs.body_y\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12925__A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13520__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19032_ net1193 _00262_ _00703_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[77\]
+ sky130_fd_sc_hd__dfrtp_1
X_16244_ net244 _02248_ net237 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__or3_4
X_13456_ net684 _07018_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__or2_1
XFILLER_0_250_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10668_ game.CPU.applesa.ab.absxs.body_x\[17\] _04699_ _04700_ game.CPU.applesa.ab.absxs.body_x\[13\]
+ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__a22o_1
XANTENNA__11549__B1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_309_Right_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16116__B net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12407_ _03240_ game.CPU.applesa.twoapples.absxs.next_head\[3\] game.CPU.applesa.twoapples.absxs.next_head\[4\]
+ _03308_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15020__B net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_341_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11013__A2 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16175_ _02181_ _02186_ _02178_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__and3b_2
X_13387_ _06872_ _06885_ net679 vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_212_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10599_ net929 game.CPU.applesa.ab.absxs.body_x\[92\] vssd1 vssd1 vccd1 vccd1 _04671_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_88_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10445__A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16488__B1 _02435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15126_ net1208 net1234 game.CPU.applesa.ab.check_walls.above.walls\[154\] vssd1
+ vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12338_ game.CPU.applesa.ab.absxs.body_y\[38\] net518 vssd1 vssd1 vccd1 vccd1 _06216_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__15955__B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10772__A1 game.CPU.applesa.ab.absxs.body_y\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19934_ clknet_leaf_42_clk game.writer.tracker.next_frame\[529\] net1327 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[529\] sky130_fd_sc_hd__dfrtp_1
X_15057_ net1212 net1238 game.CPU.applesa.ab.check_walls.above.walls\[85\] vssd1 vssd1
+ vccd1 vccd1 _00280_ sky130_fd_sc_hd__and3_1
X_12269_ net801 net419 vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_195_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_282_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14008_ net1052 _03452_ _03454_ net958 _07880_ vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_110_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19865_ clknet_leaf_20_clk game.writer.tracker.next_frame\[460\] net1310 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[460\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_207_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19216__Q game.CPU.applesa.ab.apple_possible\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11721__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18816_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[19\] _00553_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[19\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19194__CLK clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10180__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19796_ clknet_leaf_36_clk game.writer.tracker.next_frame\[391\] net1354 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[391\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_301_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16660__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15690__B net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15959_ game.CPU.applesa.ab.check_walls.above.walls\[31\] net434 vssd1 vssd1 vccd1
+ vccd1 _01971_ sky130_fd_sc_hd__nor2_1
XFILLER_0_179_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18747_ clknet_leaf_65_clk _01164_ _00484_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_179_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_223_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18059__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17204__A2 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18678_ clknet_leaf_13_clk _01095_ _00415_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[116\]
+ sky130_fd_sc_hd__dfrtp_4
X_09480_ net1091 _03476_ _03477_ net1083 vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__o22a_1
XFILLER_0_144_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17629_ game.CPU.kyle.L1.cnt_20ms\[15\] _03032_ game.CPU.kyle.L1.cnt_20ms\[16\] vssd1
+ vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a21o_1
XANTENNA__17898__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16963__A1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_349_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16176__C1 _02187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout136_A _02233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_312_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_289_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13430__S net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_288_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16026__B net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout303_A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19949__RESET_B net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17140__A1 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15865__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16313__Y _02310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16042__A game.CPU.applesa.ab.absxs.body_y\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1212_A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_257_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19537__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 net304 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_4
Xfanout312 net313 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_4
Xfanout323 game.CPU.applesa.ab.absxs.next_head\[1\] vssd1 vssd1 vccd1 vccd1 net323
+ sky130_fd_sc_hd__buf_4
Xfanout334 net335 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_4
XANTENNA_fanout672_A _07401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10515__A1 _03197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16977__A _02480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19126__Q game.CPU.applesa.ab.check_walls.above.walls\[171\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout345 game.CPU.walls.rand_wall.abduyd.next_wall\[3\] vssd1 vssd1 vccd1 vccd1
+ net345 sky130_fd_sc_hd__buf_4
XANTENNA__09381__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20005_ net1374 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
Xfanout356 _08416_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_323_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09381__B2 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ net915 game.CPU.applesa.ab.absxs.body_x\[25\] _03281_ net1107 _04056_ vssd1
+ vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__a221o_1
Xfanout367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_4
Xfanout378 net380 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_4
Xfanout389 _05864_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_161_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14257__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18965__Q game.CPU.applesa.ab.check_walls.above.walls\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09747_ net1161 game.CPU.applesa.ab.check_walls.above.walls\[68\] vssd1 vssd1 vccd1
+ vccd1 _03990_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout460_X net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18561__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19687__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_A _03190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_190_Right_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09678_ net909 game.CPU.applesa.ab.absxs.body_y\[103\] game.CPU.applesa.ab.absxs.body_y\[100\]
+ net893 vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__a22o_1
XFILLER_0_271_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11633__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16954__A1 _02408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_327_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09878__X _04121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11640_ net566 _05523_ _05524_ net746 _05528_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__a221o_1
XANTENNA__14965__B1 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__B net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12976__C1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_X clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_343_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_159_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_342_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_308_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16706__A1 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ game.CPU.applesa.ab.check_walls.above.walls\[130\] net765 vssd1 vssd1 vccd1
+ vccd1 _05460_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_172_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13310_ net483 _06748_ _07183_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__a21o_1
X_10522_ net933 game.CPU.applesa.ab.absxs.body_x\[57\] vssd1 vssd1 vccd1 vccd1 _04635_
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_250_Left_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14290_ _08158_ _08163_ vssd1 vssd1 vccd1 vccd1 _08164_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_91_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12464__B net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19067__CLK net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13615__S1 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13241_ net209 _07108_ _07114_ net284 vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__o211a_1
X_10453_ _04358_ _04586_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_268_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_296_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13172_ _07000_ _07014_ _07045_ net248 net189 vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__a221o_1
X_10384_ _03191_ game.CPU.applesa.good_collision2 _04529_ _04536_ vssd1 vssd1 vccd1
+ vccd1 _01268_ sky130_fd_sc_hd__a22o_1
XANTENNA__17131__A1 _02390_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_288_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_248_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10754__B2 game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12123_ game.CPU.applesa.ab.check_walls.above.walls\[175\] net295 net289 game.CPU.applesa.ab.check_walls.above.walls\[174\]
+ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__a22o_1
X_17980_ net590 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_264_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_263_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_261_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16931_ _02365_ _02636_ net713 vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__o21a_1
X_12054_ net816 net297 net291 game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1
+ vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__a22o_1
XFILLER_0_236_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16887__A _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19036__Q game.CPU.applesa.ab.check_walls.above.walls\[81\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18904__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ game.CPU.applesa.ab.absxs.body_y\[53\] net405 vssd1 vssd1 vccd1 vccd1 _04895_
+ sky130_fd_sc_hd__nand2_1
X_16862_ net133 _02415_ _02608_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__and3_1
X_19650_ clknet_leaf_21_clk game.writer.tracker.next_frame\[245\] net1337 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[245\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_183_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14248__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18601_ clknet_leaf_64_clk _01021_ _00338_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[82\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_125_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout890 _03368_ vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__buf_4
X_15813_ game.CPU.applesa.ab.check_walls.above.walls\[57\] net473 net468 game.CPU.applesa.ab.check_walls.above.walls\[58\]
+ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__a22o_1
X_19581_ clknet_leaf_31_clk game.writer.tracker.next_frame\[176\] net1285 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[176\] sky130_fd_sc_hd__dfrtp_4
X_16793_ _02471_ net102 _02599_ net1499 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[204\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18532_ net586 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__inv_2
XANTENNA__11824__A game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13551__S0 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15744_ net785 net450 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10809__A2 _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12956_ _06758_ _06759_ net679 vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18463_ net654 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__inv_2
X_11907_ net573 _05282_ _05283_ net750 vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_259_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ game.CPU.applesa.ab.check_walls.above.walls\[9\] net351 vssd1 vssd1 vccd1
+ vccd1 _01687_ sky130_fd_sc_hd__nand2_1
XANTENNA__15015__B net1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12887_ _06759_ _06760_ net504 vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__mux2_1
X_17414_ _02826_ _02842_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__nor2_1
X_14626_ game.CPU.clock1.counter\[13\] game.CPU.clock1.counter\[14\] _08470_ vssd1
+ vssd1 vccd1 vccd1 _08474_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_272_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11838_ net572 _05426_ _05429_ net747 vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__a22o_1
X_18394_ net619 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12967__C1 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17345_ game.CPU.kyle.L1.nextState\[1\] net1259 vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__nand2_2
XFILLER_0_157_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14557_ net1176 game.CPU.walls.rand_wall.logic_enable game.CPU.walls.abc.number_out\[4\]
+ _04256_ _08413_ vssd1 vssd1 vccd1 vccd1 _08425_ sky130_fd_sc_hd__a311oi_4
X_11769_ _03451_ net310 vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12431__B2 game.CPU.applesa.ab.absxs.body_y\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_299_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15031__A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13508_ net220 _07307_ _07381_ net284 vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_136_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17276_ net137 net113 _02336_ net733 vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__o31a_1
X_14488_ _08355_ _08356_ _08358_ _08361_ vssd1 vssd1 vccd1 vccd1 _08362_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_12_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16173__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_302_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19015_ net1196 _00244_ _00686_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_16227_ net177 net141 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__nor2_1
X_13439_ _06923_ _06926_ net702 vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10175__A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16414__X _02383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12734__A2 _06572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16158_ _01654_ _01659_ _01662_ _02102_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__o31a_1
XANTENNA__15685__B net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17122__A1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10745__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15109_ net1204 net1230 game.CPU.applesa.ab.check_walls.above.walls\[137\] vssd1
+ vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_310_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16089_ _02094_ _02095_ _02098_ _02100_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__or4_1
X_08980_ game.CPU.applesa.ab.absxs.body_x\[94\] vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_292_Right_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_283_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19917_ clknet_leaf_24_clk game.writer.tracker.next_frame\[512\] net1339 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[512\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_225_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18584__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_299_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09363__A1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__B2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19848_ clknet_leaf_40_clk game.writer.tracker.next_frame\[443\] net1356 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[443\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13790__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ net1100 game.CPU.applesa.ab.absxs.body_x\[73\] vssd1 vssd1 vccd1 vccd1 _03844_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__18785__Q game.CPU.applesa.ab.absxs.body_x\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19779_ clknet_leaf_26_clk game.writer.tracker.next_frame\[374\] net1313 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[374\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13425__S net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09532_ net1129 net811 vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__xor2_1
XANTENNA__17189__A1 _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14110__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12549__B net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ net1126 net1135 net1144 net1154 vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__or4_1
XANTENNA__16936__A1 _02369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout253_A _05210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_294_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09698__X _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09394_ _03628_ _03629_ _03633_ _03634_ _03631_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_236_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_309_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14411__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12958__C1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12422__A1 game.CPU.applesa.ab.absxs.body_x\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09858__B game.CPU.applesa.ab.absxs.body_x\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12422__B2 game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_34_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14109__X _07983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout518_A _06214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12284__B net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16324__X _02318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14780__A game.CPU.randy.counter1.count\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18252__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1048_X net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_277_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13383__C1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13922__A1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17113__A1 _02512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13922__B2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15595__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10736__A1 game.CPU.applesa.ab.absxs.body_y\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_clk_X clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_325_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10736__B2 game.CPU.applesa.ab.absxs.body_y\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18927__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout887_A _03368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09593__B game.CPU.applesa.ab.absxs.body_y\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1215_X net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14478__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_245_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1107 net1108 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__buf_4
Xfanout120 net121 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_4
Xfanout1118 game.CPU.bodymain1.main.score\[3\] vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout131 net132 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_2
XANTENNA__10532__B _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1129 game.CPU.applesa.ab.snake_head_y\[3\] vssd1 vssd1 vccd1 vccd1 net1129
+ sky130_fd_sc_hd__clkbuf_8
Xfanout142 net143 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_2
XANTENNA__09354__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout153 net155 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09354__B2 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout164 net165 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout175 net176 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_4
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_4
XFILLER_0_346_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ game.writer.tracker.frame\[368\] game.writer.tracker.frame\[369\] net1012
+ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__mux2_1
XANTENNA__13989__A1 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13790_ game.writer.tracker.frame\[429\] game.writer.tracker.frame\[431\] game.writer.tracker.frame\[432\]
+ game.writer.tracker.frame\[430\] net977 net1020 vssd1 vssd1 vccd1 vccd1 _07664_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13989__B2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_336_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ game.writer.tracker.frame\[70\] game.writer.tracker.frame\[71\] net1026 vssd1
+ vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__mux2_1
XANTENNA__16927__A1 _02359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11931__X _05819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15460_ _01440_ _01462_ _01484_ _01486_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_120_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ game.writer.updater.commands.mode\[2\] _06544_ _06546_ vssd1 vssd1 vccd1
+ vccd1 game.wr sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14411_ game.CPU.applesa.ab.absxs.body_x\[47\] net873 net961 _03310_ vssd1 vssd1
+ vccd1 vccd1 _08285_ sky130_fd_sc_hd__a22o_1
X_11623_ game.CPU.applesa.ab.check_walls.above.walls\[184\] net776 vssd1 vssd1 vccd1
+ vccd1 _05512_ sky130_fd_sc_hd__xor2_1
XFILLER_0_166_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13610__A0 game.writer.tracker.frame\[257\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15391_ _08919_ _08922_ _08926_ _08932_ vssd1 vssd1 vccd1 vccd1 _08933_ sky130_fd_sc_hd__or4b_2
XANTENNA__09768__B net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_22_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
X_17130_ _02372_ _02387_ net71 net725 vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__o31a_1
XFILLER_0_231_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14342_ game.CPU.applesa.ab.absxs.body_x\[37\] net884 net860 game.CPU.applesa.ab.absxs.body_y\[39\]
+ vssd1 vssd1 vccd1 vccd1 _08216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_181_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11554_ net775 _05442_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19702__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17061_ _02435_ net83 _02688_ net1645 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[383\]
+ sky130_fd_sc_hd__a22o_1
X_10505_ net1267 _04623_ _04624_ game.CPU.applesa.ab.absxs.body_x\[72\] vssd1 vssd1
+ vccd1 vccd1 _01187_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14273_ net1269 net883 net871 game.CPU.applesa.ab.absxs.body_y\[48\] vssd1 vssd1
+ vccd1 vccd1 _08147_ sky130_fd_sc_hd__o2bb2a_1
X_11485_ game.CPU.applesa.ab.check_walls.above.walls\[52\] net253 vssd1 vssd1 vccd1
+ vccd1 _05374_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_162_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16012_ _03238_ net344 vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__xnor2_1
X_13224_ game.writer.tracker.frame\[386\] game.writer.tracker.frame\[387\] net1038
+ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__mux2_1
XANTENNA__13913__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_347_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17104__A1 _02343_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13913__B2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10436_ game.CPU.applesa.ab.absxs.body_x\[5\] _04156_ _04159_ net1444 vssd1 vssd1
+ vccd1 vccd1 _01208_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19453__RESET_B net1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19852__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13155_ _07027_ _07028_ net514 vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_283_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10367_ game.CPU.applesa.ab.absxs.body_y\[6\] _04156_ net754 net1895 vssd1 vssd1
+ vccd1 vccd1 _01275_ sky130_fd_sc_hd__o22a_1
XANTENNA__16888__Y _02638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13126__C1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12106_ net818 net296 vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__or2_1
XANTENNA__11538__B net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13086_ game.writer.tracker.frame\[206\] game.writer.tracker.frame\[207\] net1010
+ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17963_ net656 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__inv_2
X_10298_ net1206 game.CPU.walls.rand_wall.input2 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13677__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_256_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19702_ clknet_leaf_31_clk game.writer.tracker.next_frame\[297\] net1281 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[297\] sky130_fd_sc_hd__dfrtp_1
X_16914_ _02491_ net95 _02646_ net1858 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[278\]
+ sky130_fd_sc_hd__a22o_1
X_12037_ net791 net288 net293 game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1
+ vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_251_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16410__A _02301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__A1 game.CPU.applesa.ab.absxs.body_x\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17894_ net643 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__inv_2
XFILLER_0_217_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_256_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19633_ clknet_leaf_28_clk game.writer.tracker.next_frame\[228\] net1289 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[228\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16845_ net235 net196 _02618_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__or3_2
XFILLER_0_217_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11554__A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16776_ _02436_ net64 _02594_ net1930 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[192\]
+ sky130_fd_sc_hd__a22o_1
X_19564_ clknet_leaf_34_clk game.writer.tracker.next_frame\[159\] net1329 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[159\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_189_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_220_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13988_ net1064 _03387_ _03389_ net961 _07861_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12369__B net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15727_ _03251_ net351 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__xnor2_1
X_18515_ net584 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__inv_2
XANTENNA__09024__A game.CPU.applesa.ab.absxs.body_x\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12939_ net211 _06718_ _06812_ net287 vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_17_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19495_ clknet_leaf_25_clk game.writer.tracker.next_frame\[90\] net1321 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[90\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16918__A1 _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_319_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_238_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18446_ net592 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__inv_2
X_15658_ game.CPU.applesa.ab.check_walls.above.walls\[48\] net273 vssd1 vssd1 vccd1
+ vccd1 _01670_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_14_Left_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14609_ game.CPU.clock1.counter\[7\] _08460_ game.CPU.clock1.counter\[8\] vssd1 vssd1
+ vccd1 vccd1 _08463_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18377_ net597 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15589_ game.CPU.applesa.ab.check_walls.above.walls\[35\] net461 net454 net824 _01600_
+ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_13_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17328_ net1539 _02764_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[574\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__19382__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17259_ net204 net111 net53 _02745_ net1893 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[524\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__15696__A game.CPU.applesa.ab.absxs.body_y\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_342_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10109__S _04311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_231_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13365__C1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09694__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13928__B game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__A1 game.CPU.applesa.ab.absxs.body_y\[52\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16304__B _02301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload38_A clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11288__X _05178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09536__A1_N net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14105__A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Left_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09981__X _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ net1166 vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16320__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_320_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1008_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13155__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_316_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14093__B1 game.CPU.applesa.ab.check_walls.above.walls\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12279__B net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09515_ _03756_ _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__nand2_1
XANTENNA__11183__B net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16909__A1 _02484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13840__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_X net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11300__D1 _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09446_ net914 game.CPU.applesa.ab.check_walls.above.walls\[137\] game.CPU.applesa.ab.check_walls.above.walls\[139\]
+ net925 vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_337_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19725__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13818__S1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_332_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09377_ net1150 net830 vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12295__A game.CPU.applesa.ab.check_walls.above.walls\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15593__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19964__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_331_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_312_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19875__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_305_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ _05009_ _05010_ _05012_ _05013_ _05159_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16214__B _02172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09575__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ _04408_ _04411_ _04413_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09575__B2 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14015__A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11382__B2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10152_ _04343_ _04345_ _04346_ _04344_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__o22a_2
XANTENNA__11358__B net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09327__A1 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09327__B2 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13754__S0 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10083_ _04227_ _04275_ _04229_ _04222_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__a211o_1
X_14960_ _08657_ _08666_ _08736_ vssd1 vssd1 vccd1 vccd1 _08737_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_167_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_342_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16860__A3 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout71_X net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16230__A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_233_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_293_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08948__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 game.CPU.up_button.sync1.Q vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ net1060 _03444_ net794 net852 _07781_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__a221o_1
XFILLER_0_261_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_233_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14891_ _08666_ _08667_ vssd1 vssd1 vccd1 vccd1 _08668_ sky130_fd_sc_hd__and2b_1
X_16630_ _02299_ _02518_ _02532_ net1635 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[107\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_214_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13842_ game.writer.tracker.frame\[525\] net835 net671 game.writer.tracker.frame\[528\]
+ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__o22a_1
XFILLER_0_214_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16884__B net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12189__B net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16561_ net114 net158 _02322_ net729 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__o31a_1
XANTENNA__11093__B net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13773_ game.writer.tracker.frame\[154\] net844 net712 game.writer.tracker.frame\[155\]
+ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__o22a_1
XANTENNA__13831__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ _04865_ _04869_ _04873_ _04874_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__or4_1
XFILLER_0_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15512_ _06549_ _06562_ _01505_ _01508_ _01534_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__o32a_1
X_18300_ net641 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
X_12724_ net992 net965 vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19280_ clknet_leaf_68_clk _01329_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.count\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09779__A net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16492_ net171 _02437_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_256_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_242_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18231_ net665 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
X_15443_ _08933_ _01468_ _08879_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ game.CPU.applesa.ab.absxs.body_y\[67\] net365 net525 game.CPU.applesa.ab.absxs.body_y\[65\]
+ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_182_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_178_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_328_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_316_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18162_ net589 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__inv_2
X_11606_ game.CPU.applesa.ab.check_walls.above.walls\[96\] net779 vssd1 vssd1 vccd1
+ vccd1 _05495_ sky130_fd_sc_hd__xnor2_1
X_15374_ _08898_ _08915_ vssd1 vssd1 vccd1 vccd1 _08916_ sky130_fd_sc_hd__nor2_1
XANTENNA__16128__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12586_ game.CPU.applesa.ab.absxs.body_x\[88\] net381 vssd1 vssd1 vccd1 vccd1 _06463_
+ sky130_fd_sc_hd__xnor2_2
XANTENNA__17325__B2 _02275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19984__Q game.CPU.applesa.y\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17113_ _02512_ _02692_ _02706_ net1834 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[417\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13588__X _07462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11070__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14325_ game.CPU.applesa.ab.absxs.body_y\[72\] net986 vssd1 vssd1 vccd1 vccd1 _08199_
+ sky130_fd_sc_hd__xor2_1
X_11537_ game.CPU.applesa.ab.check_walls.above.walls\[147\] net760 vssd1 vssd1 vccd1
+ vccd1 _05426_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18093_ net606 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold409 game.writer.tracker.frame\[470\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
X_17044_ _02404_ net85 _02684_ net1531 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[370\]
+ sky130_fd_sc_hd__a22o_1
X_14256_ net1267 net890 net878 game.CPU.applesa.ab.absxs.body_x\[78\] vssd1 vssd1
+ vccd1 vccd1 _08130_ sky130_fd_sc_hd__a2bb2o_1
X_11468_ net565 _05351_ _05352_ _05354_ _05355_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_40_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13207_ net512 _07078_ _07080_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10419_ game.CPU.left_button.eD1.Q1 _04563_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_267_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10453__A _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14187_ _03282_ net1046 net871 game.CPU.applesa.ab.absxs.body_y\[16\] _08060_ vssd1
+ vssd1 vccd1 vccd1 _08061_ sky130_fd_sc_hd__a221o_1
X_11399_ net746 _05283_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_209_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11373__B2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ _07008_ _07009_ _07010_ _07011_ net482 net676 vssd1 vssd1 vccd1 vccd1 _07012_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_280_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_209_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ net1195 _00222_ _00666_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[40\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13114__A2 _06985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13069_ game.writer.tracker.frame\[200\] game.writer.tracker.frame\[201\] net1015
+ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__mux2_2
XFILLER_0_188_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17946_ net628 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_2_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15795__A2_N net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_240_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11676__A2 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17877_ net636 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_355_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19616_ clknet_leaf_21_clk game.writer.tracker.next_frame\[211\] net1336 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[211\] sky130_fd_sc_hd__dfrtp_1
X_16828_ _02453_ net143 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__and2b_1
XANTENNA__16603__A3 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18622__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_356_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19748__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12099__B net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19547_ clknet_leaf_49_clk game.writer.tracker.next_frame\[142\] net1279 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[142\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13822__B1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16759_ net185 _02410_ net109 _02589_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[180\]
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_204_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12667__X game.CPU.applesa.twoapples.absxs.collision vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_278_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09300_ net1107 _03423_ _03425_ net1147 _03530_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09689__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19478_ clknet_leaf_20_clk game.writer.tracker.next_frame\[73\] net1315 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[73\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_347_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_291_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09231_ game.CPU.applesa.ab.check_walls.above.walls\[185\] vssd1 vssd1 vccd1 vccd1
+ _03480_ sky130_fd_sc_hd__inv_2
X_18429_ net586 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__inv_2
XANTENNA__11731__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18772__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19898__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_233_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09162_ game.CPU.applesa.ab.check_walls.above.walls\[57\] vssd1 vssd1 vccd1 vccd1
+ _03411_ sky130_fd_sc_hd__inv_2
XANTENNA__13050__A1 game.writer.tracker.frame\[257\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16119__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13939__A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ game.CPU.applesa.ab.absxs.body_y\[48\] vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout216_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19128__CLK net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_309_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16034__B net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__B net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09557__A1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09557__B2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1125_A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16827__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15873__B net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11178__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ game.CPU.apple_location\[4\] game.CPU.applesa.ab.apple_location\[4\] _04207_
+ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__mux2_1
XANTENNA__19278__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout585_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09309__A1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09309__B2 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ net1116 vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__inv_2
XFILLER_0_283_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16050__A game.CPU.applesa.ab.absxs.body_y\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12313__B1 _06163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13510__C1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10810__B _04702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19134__Q game.CPU.applesa.ab.check_walls.above.walls\[179\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout540_X net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17004__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_333_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10770_ game.CPU.applesa.ab.absxs.body_y\[74\] _04675_ _04676_ game.CPU.applesa.ab.absxs.body_y\[70\]
+ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__a22o_1
X_09429_ game.CPU.applesa.ab.snake_head_x\[2\] _03440_ _03668_ _03669_ _03670_ vssd1
+ vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__a221o_1
XFILLER_0_176_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12440_ game.CPU.applesa.ab.absxs.body_x\[104\] net382 vssd1 vssd1 vccd1 vccd1 _06317_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_191_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09886__X _04129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13041__A1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10257__B net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09796__A1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ game.CPU.applesa.ab.absxs.body_x\[115\] net530 vssd1 vssd1 vccd1 vccd1 _06248_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09796__B2 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16225__A net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14110_ net938 game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1 vssd1 vccd1
+ vccd1 _07984_ sky130_fd_sc_hd__xor2_1
X_11322_ game.CPU.applesa.ab.check_walls.above.walls\[68\] net253 vssd1 vssd1 vccd1
+ vccd1 _05211_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_278_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15090_ net1211 net1237 net797 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__and3_1
XFILLER_0_278_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_344_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14041_ net877 game.CPU.applesa.ab.check_walls.above.walls\[114\] game.CPU.applesa.ab.check_walls.above.walls\[115\]
+ net876 _07914_ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__o221a_1
XANTENNA__11369__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11253_ _05128_ _05129_ _05131_ _05133_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__or4_1
X_10204_ net1089 _04394_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__nor2_1
XANTENNA__11088__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15783__B net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17086__A3 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ _03234_ net416 vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__nand2_1
XANTENNA__16294__A1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08949__Y _03199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17800_ net1049 _03134_ _03139_ _01548_ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__o211a_1
XANTENNA__13727__S0 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ game.CPU.randy.f1.c1.count\[10\] game.CPU.randy.f1.c1.count\[13\] game.CPU.randy.f1.c1.count\[12\]
+ game.CPU.randy.f1.c1.count\[15\] vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__or4_1
X_18780_ clknet_leaf_64_clk _01197_ _00517_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_15992_ _03435_ game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 _02004_ sky130_fd_sc_hd__nor2_1
XANTENNA__18645__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14399__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13501__C1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ _04239_ _04273_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__nor2_1
X_17731_ _03085_ _03096_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__nor2_1
X_14943_ _08714_ _08717_ _08719_ vssd1 vssd1 vccd1 vccd1 _08720_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12855__A1 game.writer.tracker.frame\[305\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11658__A2 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13871__X _07745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17343__X _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17662_ _08811_ _03009_ _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__or3_1
X_14874_ game.CPU.walls.abc.number\[6\] game.CPU.walls.abc.number\[2\] game.CPU.walls.abc.counter
+ vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__mux2_1
XANTENNA__15007__C game.CPU.applesa.ab.check_walls.above.walls\[35\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_230_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19401_ clknet_leaf_47_clk _01401_ net1279 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.x\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_13825_ net178 _07638_ _07660_ _07698_ net191 vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__a311o_1
X_16613_ game.writer.tracker.frame\[101\] _02515_ vssd1 vssd1 vccd1 vccd1 _02523_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_214_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17593_ _03001_ _03011_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__or2_1
XANTENNA__18795__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13804__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16544_ net202 net146 _02393_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__and3_1
X_19332_ clknet_leaf_72_clk net1429 _00937_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twomode.number\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13756_ _07628_ _07629_ net482 vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__mux2_1
X_10968_ _03227_ net319 vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_329_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12707_ _06554_ _06564_ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__xor2_1
XANTENNA__11551__B net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16475_ _02274_ _02425_ net737 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19263_ clknet_leaf_9_clk _00051_ _00893_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_13687_ _07559_ _07560_ net477 vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__mux2_1
X_10899_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__inv_2
X_15426_ game.writer.updater.commands.cmd_num\[0\] _08934_ _01453_ vssd1 vssd1 vccd1
+ vccd1 _01454_ sky130_fd_sc_hd__o21a_2
X_18214_ net666 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__inv_2
XANTENNA__13032__A1 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19194_ clknet_leaf_46_clk net338 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.y_final\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12638_ _06323_ _06467_ _06325_ _06466_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__or4b_2
XFILLER_0_155_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15958__B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10167__B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16406__Y _02376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15357_ _08885_ _08898_ vssd1 vssd1 vccd1 vccd1 _08899_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18145_ net630 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__inv_2
X_12569_ game.CPU.applesa.ab.absxs.body_x\[117\] net378 net520 game.CPU.applesa.ab.absxs.body_y\[118\]
+ _06445_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__o221a_1
XANTENNA__13111__X _06985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_215_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11594__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14308_ _03248_ net1061 net876 game.CPU.applesa.ab.absxs.body_x\[31\] _08178_ vssd1
+ vssd1 vccd1 vccd1 _08182_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18076_ net658 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__inv_2
Xwire181 _06638_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_2
Xhold206 game.writer.tracker.frame\[366\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
X_15288_ _08814_ _08832_ vssd1 vssd1 vccd1 vccd1 _08839_ sky130_fd_sc_hd__nor2_1
Xhold217 game.writer.tracker.frame\[447\] vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xwire192 _05720_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12382__B net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_300_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold228 game.writer.tracker.frame\[109\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
X_17027_ _02524_ _02663_ _02680_ net1821 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[357\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09539__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19420__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 game.writer.tracker.frame\[166\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ game.CPU.applesa.ab.absxs.body_y\[114\] net953 vssd1 vssd1 vccd1 vccd1 _08113_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__09539__B2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10183__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_278_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16422__X _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout708 net709 vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_4
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15693__B net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout719 net726 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_41_clk_X clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13718__S0 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16285__B2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ net1127 net789 vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__or2_1
XFILLER_0_265_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18978_ net1199 _00203_ _00649_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19570__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17929_ net659 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__inv_2
XANTENNA__10630__B game.CPU.applesa.ab.absxs.body_x\[53\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14102__B net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1290 net1293 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13941__B game.CPU.applesa.ab.check_walls.above.walls\[66\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15796__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_354_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19556__RESET_B net1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09212__A game.CPU.applesa.ab.check_walls.above.walls\[157\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11461__B net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout333_A game.CPU.walls.rand_wall.abduyd.next_wall\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1075_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09214_ net788 vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_315_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14220__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16760__A2 _02412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13669__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1 vccd1 vccd1
+ _03394_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout121_X net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout500_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1242_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout219_X net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09076_ game.CPU.applesa.ab.absxs.body_y\[97\] vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__inv_2
XANTENNA__16512__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19129__Q game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12292__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15884__A game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18260__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18668__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1128_X net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19913__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_338_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout967_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13709__S0 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13608__S net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ net1158 net1262 vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__or2_1
XFILLER_0_338_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14287__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout79_A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_164_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_354_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09702__A1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ net787 net300 vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__nand2_1
XANTENNA__09702__B2 net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_354_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17240__A3 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ game.CPU.applesa.ab.check_walls.above.walls\[5\] net309 vssd1 vssd1 vccd1
+ vccd1 _05759_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13610_ game.writer.tracker.frame\[257\] game.writer.tracker.frame\[259\] game.writer.tracker.frame\[260\]
+ game.writer.tracker.frame\[258\] net967 net996 vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__mux4_1
XFILLER_0_196_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10822_ net1443 game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__nor2_2
X_14590_ net739 net331 vssd1 vssd1 vccd1 vccd1 _08452_ sky130_fd_sc_hd__nor2_1
XFILLER_0_357_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09466__B1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12467__B net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13541_ game.writer.tracker.frame\[113\] game.writer.tracker.frame\[115\] game.writer.tracker.frame\[116\]
+ game.writer.tracker.frame\[114\] net978 net1015 vssd1 vssd1 vccd1 vccd1 _07415_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_253_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10753_ game.CPU.applesa.ab.absxs.body_y\[110\] _04665_ _04666_ game.CPU.applesa.ab.absxs.body_y\[106\]
+ vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11812__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16260_ net248 _02265_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__or2_2
XFILLER_0_82_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13472_ _07074_ _07075_ net704 vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_299_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15778__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10684_ game.CPU.applesa.ab.absxs.body_x\[8\] _04689_ _04707_ game.CPU.applesa.ab.absxs.body_x\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__a22o_1
XFILLER_0_326_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16751__A2 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ game.CPU.applesa.normal1.number\[3\] _08773_ vssd1 vssd1 vccd1 vccd1 _08778_
+ sky130_fd_sc_hd__or2_1
X_12423_ game.CPU.applesa.ab.absxs.body_y\[33\] net523 net363 game.CPU.applesa.ab.absxs.body_y\[32\]
+ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_117_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19443__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16191_ _02126_ _02129_ _02201_ _02202_ _01793_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__o41a_1
XFILLER_0_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15142_ net1209 net1235 game.CPU.applesa.ab.check_walls.above.walls\[170\] vssd1
+ vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__and3_1
X_12354_ game.CPU.applesa.ab.absxs.body_x\[78\] net371 vssd1 vssd1 vccd1 vccd1 _06231_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_294_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13317__A2 _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ net563 _05193_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__nor2_4
X_19950_ clknet_leaf_38_clk game.writer.tracker.next_frame\[545\] net1326 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[545\] sky130_fd_sc_hd__dfrtp_1
X_15073_ net1212 net1238 net804 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12285_ _03451_ net421 vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__nor2_1
XANTENNA__19593__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18901_ clknet_leaf_69_clk _01268_ _00585_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.good_collision2
+ sky130_fd_sc_hd__dfrtp_1
X_14024_ net1052 _03466_ net786 net856 vssd1 vssd1 vccd1 vccd1 _07898_ sky130_fd_sc_hd__a22o_1
XANTENNA__09792__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11236_ _05122_ _05123_ _05124_ _05125_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_56_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19881_ clknet_leaf_26_clk game.writer.tracker.next_frame\[476\] net1319 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[476\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_264_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_248_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11879__A2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13518__S net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18832_ clknet_leaf_0_clk _01223_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_11167_ _05047_ _05050_ _05051_ _05056_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__or4_1
XFILLER_0_248_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_186_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10118_ game.CPU.applesa.enable_in game.CPU.applesa.twoapples.x_final\[1\] _03212_
+ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__a21o_1
X_18763_ clknet_leaf_51_clk _01180_ _00500_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[61\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11546__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15018__B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11098_ game.CPU.applesa.ab.absxs.body_x\[57\] net413 vssd1 vssd1 vccd1 vccd1 _04988_
+ sky130_fd_sc_hd__xnor2_1
X_15975_ _01979_ _01980_ _01984_ _01985_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a22o_1
XANTENNA__17216__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17714_ _03085_ _03086_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__nor2_1
X_14926_ _08678_ _08681_ _08683_ _08679_ _08662_ vssd1 vssd1 vccd1 vccd1 _08703_ sky130_fd_sc_hd__o311a_1
X_10049_ net1271 net846 vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__or2_4
X_18694_ clknet_leaf_59_clk _01111_ _00431_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[40\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11500__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_264_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11500__B2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17645_ _08804_ _03037_ _03042_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__and3b_1
XFILLER_0_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_353_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14857_ game.CPU.randy.f1.c1.count\[12\] _08647_ vssd1 vssd1 vccd1 vccd1 _08649_
+ sky130_fd_sc_hd__and2_1
XANTENNA__19502__Q game.writer.tracker.frame\[97\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_230_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ game.writer.tracker.frame\[445\] game.writer.tracker.frame\[447\] game.writer.tracker.frame\[448\]
+ game.writer.tracker.frame\[446\] net980 net1038 vssd1 vssd1 vccd1 vccd1 _07682_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_201_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14788_ _08605_ _08606_ net139 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_67_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17576_ net1446 net264 _02880_ _02999_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_275_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16990__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19315_ net1165 _00029_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twomode.counter
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11264__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13739_ _07611_ _07612_ net491 vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__mux2_1
X_16527_ net2056 _02463_ _02465_ net125 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[72\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_217_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_318_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19246_ clknet_leaf_17_clk _00060_ _00884_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_16458_ net240 _02367_ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__nor2_8
XANTENNA__15688__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13556__A2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15409_ _01436_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__inv_2
X_16389_ net135 net115 _02364_ _02361_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[35\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19177_ clknet_leaf_6_clk _01296_ _00839_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_332_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18128_ net578 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__inv_2
XFILLER_0_289_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_300_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10117__S _04311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18059_ net634 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11319__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_286_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10790__A2 game.CPU.applesa.ab.absxs.body_y\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09901_ _03593_ _03598_ _03694_ _03981_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkload20_A clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16258__A1 _06571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout505 net516 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_228_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout516 _06595_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_2
X_20021_ net1276 vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_09832_ _04067_ _04071_ _04072_ _04074_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__or4_2
XANTENNA__18960__CLK net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout527 _06213_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_272_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout538 net540 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14269__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_238_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout549 net550 vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_265_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09763_ net1091 game.CPU.applesa.ab.check_walls.above.walls\[98\] vssd1 vssd1 vccd1
+ vccd1 _04006_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout283_A net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19316__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09694_ net1139 game.CPU.applesa.ab.absxs.body_y\[6\] vssd1 vssd1 vccd1 vccd1 _03937_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__09696__B1 game.CPU.applesa.ab.absxs.body_y\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17222__A3 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout450_A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_317_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout169_X net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16430__A1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1192_A game.CPU.walls.rand_wall.good_spot vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_324_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_36_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16981__A2 _02460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_239_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11255__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13795__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout715_A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12855__X _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout336_X net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1078_X net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15598__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_340_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09596__B game.CPU.applesa.ab.absxs.body_y\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_161_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11558__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_350_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09128_ net954 vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_350_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09620__B1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16497__A1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14007__B game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_328_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09059_ game.CPU.applesa.ab.absxs.body_y\[52\] vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16503__A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12070_ _05955_ _05956_ _05953_ _05954_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__and4b_1
XANTENNA__18698__Q game.CPU.applesa.ab.absxs.body_x\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold570 game.CPU.applesa.ab.count\[1\] vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10822__Y _00039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold581 game.CPU.applesa.ab.absxs.body_x\[2\] vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 game.writer.tracker.frame\[453\] vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13338__S net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11021_ game.CPU.applesa.ab.absxs.body_y\[91\] net396 vssd1 vssd1 vccd1 vccd1 _04911_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__11647__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11263__A2_N net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11366__B net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15760_ game.CPU.applesa.ab.absxs.body_y\[119\] net435 vssd1 vssd1 vccd1 vccd1 _01772_
+ sky130_fd_sc_hd__xnor2_1
X_12972_ net227 _06653_ _06845_ net278 vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_51_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14310__X _08184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13483__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14711_ _03513_ _08547_ vssd1 vssd1 vccd1 vccd1 _08548_ sky130_fd_sc_hd__nand2_1
X_11923_ net782 net391 vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_339_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17213__A3 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15691_ game.CPU.applesa.ab.absxs.body_y\[31\] net431 vssd1 vssd1 vccd1 vccd1 _01703_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_200_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14642_ game.CPU.clock1.counter\[19\] game.CPU.clock1.counter\[20\] _08480_ vssd1
+ vssd1 vccd1 vccd1 _08484_ sky130_fd_sc_hd__and3_1
X_17430_ net1275 _02825_ net427 vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__and3_1
XFILLER_0_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11854_ net803 net303 net394 game.CPU.applesa.ab.check_walls.above.walls\[100\] vssd1
+ vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_157_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_318_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16972__A2 _02638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12197__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14432__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10805_ game.CPU.applesa.ab.absxs.body_y\[24\] _04695_ _04698_ game.CPU.applesa.ab.absxs.body_y\[20\]
+ vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__a22o_1
XANTENNA__11246__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13330__S1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14573_ game.CPU.clock1.counter\[3\] game.CPU.clock1.counter\[2\] game.CPU.clock1.counter\[4\]
+ game.CPU.clock1.counter\[7\] vssd1 vssd1 vccd1 vccd1 _08435_ sky130_fd_sc_hd__or4b_1
X_17361_ net1114 net1115 game.CPU.bodymain1.main.score\[7\] vssd1 vssd1 vccd1 vccd1
+ _02791_ sky130_fd_sc_hd__nor3b_2
XANTENNA__15789__A game.CPU.applesa.ab.absxs.body_y\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_345_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12765__X _06639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11785_ net822 net304 vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19100_ net1180 _00138_ _00771_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[145\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13524_ net178 _07386_ _07397_ net173 vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__a211o_2
X_16312_ _02298_ _02308_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__nor2_4
XANTENNA__11797__B2 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17292_ net183 net116 _02521_ _02753_ net1628 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[548\]
+ sky130_fd_sc_hd__a32o_1
X_10736_ game.CPU.applesa.ab.absxs.body_y\[15\] _04653_ _04654_ game.CPU.applesa.ab.absxs.body_y\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__a22o_1
XANTENNA__16185__B1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19959__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16243_ net275 _02226_ _02227_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__o21a_1
X_19031_ net1193 _00261_ _00702_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[76\]
+ sky130_fd_sc_hd__dfrtp_4
X_13455_ net705 _06996_ _07328_ net498 vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__o211a_1
XFILLER_0_353_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ game.CPU.applesa.ab.absxs.body_x\[18\] _04699_ _04700_ game.CPU.applesa.ab.absxs.body_x\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_273_Right_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_max_cap179_A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11549__B2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12406_ _06280_ _06281_ _06282_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__and3_1
X_16174_ _01623_ _02182_ _02183_ _02185_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__or4_1
X_13386_ _07258_ _07259_ net485 vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__mux2_1
XANTENNA__15020__C game.CPU.applesa.ab.check_walls.above.walls\[48\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_212_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10598_ game.CPU.applesa.ab.absxs.body_x\[97\] net263 _04670_ net929 vssd1 vssd1
+ vccd1 vccd1 _01140_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_188_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15125_ net1208 net1233 game.CPU.applesa.ab.check_walls.above.walls\[153\] vssd1
+ vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__and3_1
XFILLER_0_140_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16488__B2 _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12337_ net364 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.absxs.next_head\[7\]
+ sky130_fd_sc_hd__clkinv_4
XANTENNA__16413__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12941__A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10772__A2 _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19933_ clknet_leaf_48_clk game.writer.tracker.next_frame\[528\] net1307 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[528\] sky130_fd_sc_hd__dfrtp_1
X_15056_ net1212 net1242 net810 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__and3_1
X_12268_ net801 net419 vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__and2_1
XFILLER_0_294_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14007_ net938 game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1 vssd1 vccd1
+ vccd1 _07881_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11219_ game.CPU.applesa.ab.absxs.body_x\[37\] net321 vssd1 vssd1 vccd1 vccd1 _05109_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__15029__A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19864_ clknet_leaf_20_clk game.writer.tracker.next_frame\[459\] net1310 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[459\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_110_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10461__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19339__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ _05997_ _06084_ _05999_ _05998_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__or4bb_1
XANTENNA__11721__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_275_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18815_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[18\] _00552_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[18\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09027__A game.CPU.applesa.ab.absxs.body_x\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_207_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15971__B net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19795_ clknet_leaf_35_clk game.writer.tracker.next_frame\[390\] net1354 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[390\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15999__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16660__A1 _02243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_268_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18746_ clknet_leaf_61_clk _01163_ _00483_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_15958_ _03392_ net348 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09678__B1 game.CPU.applesa.ab.absxs.body_y\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_223_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17204__A3 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14909_ net1171 _08426_ _08428_ net1170 _08685_ vssd1 vssd1 vccd1 vccd1 _08686_ sky130_fd_sc_hd__a221o_1
XANTENNA__19489__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18677_ clknet_leaf_8_clk _01094_ _00414_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_15889_ game.CPU.applesa.ab.check_walls.above.walls\[137\] net472 vssd1 vssd1 vccd1
+ vccd1 _01901_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_203_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17628_ net2010 _03032_ _03033_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__o21a_1
XANTENNA__14423__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17559_ _02932_ _02980_ _02983_ _02984_ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__or4_1
XANTENNA__18075__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload68_A clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_312_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19229_ clknet_leaf_57_clk net1414 _00867_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.normal1.number\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_288_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_240_Right_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_258_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17140__A2 _02410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_257_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10763__A2 _04590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16042__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout498_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_319_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout313 _05600_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_4
Xfanout324 game.CPU.applesa.ab.absxs.next_head\[0\] vssd1 vssd1 vccd1 vccd1 net324
+ sky130_fd_sc_hd__clkbuf_8
Xfanout335 game.CPU.walls.rand_wall.abduyd.next_wall\[6\] vssd1 vssd1 vccd1 vccd1
+ net335 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1205_A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10515__A2 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout346 net347 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_4
XANTENNA__16977__B _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20004_ clknet_leaf_45_clk game.writer.updater.update.next\[2\] net1300 vssd1 vssd1
+ vccd1 vccd1 game.writer.updater.commands.mode\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_226_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09815_ net1136 _03349_ game.CPU.applesa.ab.absxs.body_y\[25\] net901 _04057_ vssd1
+ vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__a221o_1
XANTENNA_input3_A gpio_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_323_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15881__B net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11186__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12997__S net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 _06215_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_4
XANTENNA__18706__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout379 net380 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_2
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_253_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout665_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16651__A1 _02415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ net926 game.CPU.applesa.ab.check_walls.above.walls\[67\] _03419_ net1150
+ _03982_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__a221o_1
XFILLER_0_213_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09677_ net1093 game.CPU.applesa.ab.absxs.body_x\[102\] vssd1 vssd1 vccd1 vccd1 _03920_
+ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12298__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1195_X net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16403__B2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15105__C net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14414__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18981__Q game.CPU.applesa.ab.check_walls.above.walls\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13768__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13312__S1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11779__A1 net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_159_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_308_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11570_ game.CPU.applesa.ab.check_walls.above.walls\[131\] net759 vssd1 vssd1 vccd1
+ vccd1 _05459_ sky130_fd_sc_hd__xnor2_2
XANTENNA__16167__B1 game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16217__B net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10521_ _04634_ game.CPU.applesa.ab.absxs.body_x\[62\] net425 vssd1 vssd1 vccd1 vccd1
+ _01181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12728__A0 game.writer.tracker.frame\[98\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13240_ net226 _07113_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10452_ _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__inv_2
XANTENNA__16504__Y _02449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ net285 _07022_ _07030_ _07043_ _07044_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__o32a_1
X_10383_ net1134 _03204_ _04533_ _04534_ _04535_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__o2111a_1
XANTENNA__17131__A2 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16233__A net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10754__A2 _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_248_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12122_ _06006_ _06007_ _06008_ _06005_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__a211o_1
XANTENNA__16890__A1 _02267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11377__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_261_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16930_ _02514_ net92 _02650_ net1568 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[290\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_53_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12053_ net816 net297 net291 game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1
+ vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__o22ai_1
XANTENNA__16887__B _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ _04882_ _04889_ _04890_ _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__or4_1
XANTENNA__11096__B net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16861_ net158 _02413_ net99 net730 vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__o31a_1
XFILLER_0_263_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_183_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19631__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_244_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout880 _03372_ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_8
X_18600_ clknet_leaf_64_clk _01020_ _00337_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[81\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_69_Left_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout891 net892 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_125_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15812_ _03411_ net351 net349 _03412_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__a22o_1
X_19580_ clknet_leaf_32_clk game.writer.tracker.next_frame\[175\] net1284 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[175\] sky130_fd_sc_hd__dfrtp_1
X_16792_ _02468_ net100 net716 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__o21a_1
Xclkbuf_3_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_clk sky130_fd_sc_hd__clkbuf_8
X_18531_ net601 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__inv_2
X_12955_ net483 _06828_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__or2_1
X_15743_ _03471_ net346 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11824__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13551__S1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12664__C1 _06336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17198__A2 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14200__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_342_Right_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11906_ game.CPU.applesa.ab.check_walls.above.walls\[95\] net312 vssd1 vssd1 vccd1
+ vccd1 _05794_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_319_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18462_ net654 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12886_ game.writer.tracker.frame\[14\] game.writer.tracker.frame\[15\] net1004 vssd1
+ vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__mux2_1
X_15674_ game.CPU.applesa.ab.check_walls.above.walls\[12\] net453 vssd1 vssd1 vccd1
+ vccd1 _01686_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12001__A game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19781__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_259_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16945__A2 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17413_ _02842_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13759__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11837_ net571 _05426_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__nor2_1
X_14625_ game.CPU.clock1.counter\[13\] game.CPU.clock1.counter\[12\] _08469_ game.CPU.clock1.counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _08473_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_64_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_272_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18393_ net617 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__inv_2
XANTENNA__12936__A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12967__B1 _06840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14556_ game.CPU.walls.abc.enable game.CPU.walls.abc.number_out\[4\] vssd1 vssd1
+ vccd1 vccd1 _08424_ sky130_fd_sc_hd__nand2_1
X_17344_ _03218_ _03219_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__nor2_1
XANTENNA__16158__B1 _02102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11768_ net793 net390 net305 net792 vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_194_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12431__A2 game.CPU.applesa.twoapples.absxs.next_head\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Left_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19011__CLK net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13507_ net478 _07304_ _07306_ net202 vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__a211o_1
XANTENNA__15031__B net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ game.CPU.applesa.ab.absxs.body_y\[47\] _04640_ _04641_ game.CPU.applesa.ab.absxs.body_y\[43\]
+ vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__a22o_1
X_17275_ _02278_ _02497_ _02749_ net1890 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[536\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14487_ _08053_ _08240_ _08359_ _08360_ vssd1 vssd1 vccd1 vccd1 _08361_ sky130_fd_sc_hd__and4_1
X_11699_ net742 _05587_ _05585_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10456__A _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19014_ net1202 _00242_ _00685_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[59\]
+ sky130_fd_sc_hd__dfrtp_4
X_13438_ _07310_ _07311_ net212 vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__mux2_1
X_16226_ net175 net141 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__or2_2
XANTENNA__15966__B net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_286_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16157_ _01647_ _01649_ _01652_ _01653_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__or4_1
XFILLER_0_106_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13369_ _06686_ _06697_ net678 vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17122__A2 _02373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11942__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19161__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10745__A2 game.CPU.applesa.ab.absxs.body_y\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15108_ net1207 net1230 game.CPU.applesa.ab.check_walls.above.walls\[136\] vssd1
+ vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16088_ game.CPU.applesa.ab.check_walls.above.walls\[145\] net472 net459 game.CPU.applesa.ab.check_walls.above.walls\[147\]
+ _02099_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a221o_1
XANTENNA__12390__B game.CPU.applesa.twoapples.absxs.next_head\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_283_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18729__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19916_ clknet_leaf_24_clk game.writer.tracker.next_frame\[511\] net1339 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[511\] sky130_fd_sc_hd__dfrtp_1
X_15039_ net1219 net1244 game.CPU.applesa.ab.check_walls.above.walls\[67\] vssd1 vssd1
+ vccd1 vccd1 _00260_ sky130_fd_sc_hd__and3_1
XANTENNA__10191__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13695__A1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_225_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09899__B1 _03784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_299_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_87_Left_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19847_ clknet_leaf_40_clk game.writer.tracker.next_frame\[442\] net1355 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[442\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_242_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16633__A1 _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09600_ net926 game.CPU.applesa.ab.absxs.body_x\[75\] game.CPU.applesa.ab.absxs.body_y\[73\]
+ net900 vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_208_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19778_ clknet_leaf_26_clk game.writer.tracker.next_frame\[373\] net1312 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[373\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18879__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09531_ _03764_ _03765_ _03768_ _03773_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__or4_4
X_18729_ clknet_leaf_13_clk _01146_ _00466_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[111\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14110__B game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09462_ net1081 net1090 net1097 net1106 vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__or4_1
XFILLER_0_305_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16397__B1 _02369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_176_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16936__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_294_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09393_ net1099 _03465_ game.CPU.applesa.ab.check_walls.above.walls\[162\] net920
+ _03627_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout246_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_236_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_96_Left_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12422__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12565__B net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11630__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout413_A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1155_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19504__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14175__A2 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14780__B _04486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout201_X net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10653__X _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12581__A game.CPU.applesa.ab.absxs.body_y\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17113__A2 _02692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1322_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_325_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10736__A2 _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19137__Q game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19654__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_247_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11197__A game.CPU.applesa.ab.absxs.body_x\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15892__A game.CPU.applesa.ab.absxs.body_x\[40\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout110 _02558_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_4
Xfanout1108 net1113 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1110_X net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout121 _02633_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_245_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1119 game.CPU.bodymain1.main.score\[2\] vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__clkbuf_4
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_4
Xfanout143 _02608_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_2
XANTENNA__18976__Q game.CPU.applesa.ab.check_walls.above.walls\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
XFILLER_0_245_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout570_X net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout165 net166 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16500__B _02444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 _06700_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout187 _06589_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_4
Xfanout198 net199 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_346_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout61_A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14301__A game.CPU.applesa.ab.absxs.body_y\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09729_ net1083 game.CPU.applesa.ab.absxs.body_x\[35\] vssd1 vssd1 vccd1 vccd1 _03972_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__12646__C1 _06522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12740_ net508 _06611_ _06613_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__a21o_1
XFILLER_0_198_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09889__X _04132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_336_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16927__A2 _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19034__CLK net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12671_ game.writer.updater.commands.mode\[2\] _06545_ vssd1 vssd1 vccd1 vccd1 _06546_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_120_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16228__A net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14410_ _08280_ _08283_ _08281_ _08282_ vssd1 vssd1 vccd1 vccd1 _08284_ sky130_fd_sc_hd__or4b_1
XFILLER_0_343_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15132__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11622_ net776 _05510_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__xnor2_1
X_15390_ _08900_ _08914_ _08916_ _08931_ _08930_ vssd1 vssd1 vccd1 vccd1 _08932_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09814__B1 game.CPU.applesa.ab.absxs.body_y\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_343_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12475__B net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09130__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14341_ game.CPU.applesa.ab.absxs.body_x\[36\] net890 net963 _03312_ vssd1 vssd1
+ vccd1 vccd1 _08215_ sky130_fd_sc_hd__a22o_1
X_11553_ game.CPU.applesa.ab.check_walls.above.walls\[193\] net770 vssd1 vssd1 vccd1
+ vccd1 _05442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10276__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18443__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19184__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17060_ _02431_ net83 _02688_ net1684 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[382\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ game.CPU.applesa.ab.absxs.body_x\[77\] _04623_ _04624_ game.CPU.applesa.ab.absxs.body_x\[73\]
+ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__a22o_1
X_14272_ _08142_ _08143_ _08145_ vssd1 vssd1 vccd1 vccd1 _08146_ sky130_fd_sc_hd__or3b_1
XANTENNA__16560__B1 _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11484_ _03409_ net317 vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15786__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16011_ net1270 net434 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__xnor2_1
X_13223_ game.writer.tracker.frame\[390\] game.writer.tracker.frame\[391\] net1039
+ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12177__B2 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10435_ game.CPU.applesa.ab.absxs.body_x\[6\] net847 _04158_ net1966 vssd1 vssd1
+ vccd1 vccd1 _01209_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_347_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17104__A2 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13154_ game.writer.tracker.frame\[182\] game.writer.tracker.frame\[183\] net1036
+ vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__mux2_1
X_10366_ game.CPU.applesa.ab.absxs.body_y\[7\] net850 _04158_ net1453 vssd1 vssd1
+ vccd1 vccd1 _01276_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_131_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19047__Q game.CPU.applesa.ab.check_walls.above.walls\[92\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12105_ net797 net292 net295 game.CPU.applesa.ab.check_walls.above.walls\[119\] vssd1
+ vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__o2bb2a_1
X_13085_ net502 _06956_ _06958_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__a21o_1
X_17962_ net657 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__inv_2
X_10297_ _03214_ net1441 _04473_ _04481_ vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__o31a_1
X_19701_ clknet_leaf_30_clk game.writer.tracker.next_frame\[296\] net1284 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[296\] sky130_fd_sc_hd__dfrtp_1
X_16913_ _02489_ net95 _02646_ net1767 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[277\]
+ sky130_fd_sc_hd__a22o_1
X_12036_ _05920_ _05921_ _05922_ _05919_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a211o_1
XFILLER_0_252_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_256_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17893_ net620 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__inv_2
XANTENNA__19422__RESET_B net1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__A2 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19632_ clknet_leaf_27_clk game.writer.tracker.next_frame\[227\] net1309 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[227\] sky130_fd_sc_hd__dfrtp_1
X_16844_ net971 _02246_ _02305_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13429__A1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_256_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09305__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19563_ clknet_leaf_37_clk game.writer.tracker.next_frame\[158\] net1329 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[158\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15026__B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16775_ _02432_ _02561_ net736 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__o21a_1
X_13987_ net1073 _03386_ _03388_ net1059 vssd1 vssd1 vccd1 vccd1 _07861_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_358_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18514_ net579 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__inv_2
X_15726_ _03240_ net344 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17522__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12938_ net493 _06811_ _06810_ net228 vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__o211a_1
X_19494_ clknet_leaf_24_clk game.writer.tracker.next_frame\[89\] net1338 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[89\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12652__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_272_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17040__A1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18445_ net592 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__inv_2
XANTENNA__10663__B2 game.CPU.applesa.ab.absxs.body_x\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15657_ _03409_ net339 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__xnor2_1
X_12869_ game.writer.tracker.frame\[294\] game.writer.tracker.frame\[295\] net988
+ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14608_ net1492 _08460_ _08462_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[7\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19527__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18376_ net597 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__inv_2
X_15588_ net822 net440 net474 game.CPU.applesa.ab.check_walls.above.walls\[33\] vssd1
+ vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_306_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12385__B net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17327_ net1722 _02764_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[573\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_7_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14539_ game.writer.control.current\[0\] game.writer.control.current\[1\] _06547_
+ vssd1 vssd1 vccd1 vccd1 _08412_ sky130_fd_sc_hd__and3b_1
XANTENNA__14881__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_300_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17258_ _02275_ _02300_ _02745_ net1813 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[523\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15696__B net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16551__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_231_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18551__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19677__CLK clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16209_ _02019_ _02022_ _02023_ _02220_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__or4_2
XFILLER_0_302_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09694__B game.CPU.applesa.ab.absxs.body_y\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17189_ _02496_ net78 _02728_ net1721 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[471\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_287_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10718__A2 _04609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_297_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14105__B game.CPU.applesa.ab.check_walls.above.walls\[49\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08962_ game.CPU.applesa.twoapples.start_enable vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__inv_2
XFILLER_0_227_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16160__X _02172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17416__B _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16320__B net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout196_A _02289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13436__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_320_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_242_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_242_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11464__B net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14093__A1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14093__B2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ net1085 _03271_ game.CPU.applesa.ab.absxs.body_x\[48\] net912 vssd1 vssd1
+ vccd1 vccd1 _03757_ sky130_fd_sc_hd__o22a_1
XANTENNA__13960__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11300__C1 _05185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17031__A1 _02375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ net1106 game.CPU.applesa.ab.check_walls.above.walls\[136\] vssd1 vssd1 vccd1
+ vccd1 _03688_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout151_X net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout530_A net532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1272_A net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14494__C _08366_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11480__A game.CPU.applesa.ab.check_walls.above.walls\[48\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_332_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09376_ net1094 game.CPU.applesa.ab.check_walls.above.walls\[10\] vssd1 vssd1 vccd1
+ vccd1 _03619_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15593__B2 game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12295__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15887__A game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_331_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1060_X net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18263__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1158_X net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_340_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09885__A _04121_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout997_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_320_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17098__A1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19933__RESET_B net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ _04373_ _04388_ _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__nor3_1
XANTENNA__16214__C _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11639__B net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13108__B1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15648__A2 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10151_ net1260 game.CPU.randy.f1.state\[3\] game.CPU.randy.f1.state\[2\] vssd1 vssd1
+ vccd1 vccd1 _04346_ sky130_fd_sc_hd__or3b_1
XANTENNA__13203__S0 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14320__A2 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10082_ _04221_ _04289_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_167_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_342_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout952_X net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ _07777_ _07778_ _07779_ _07780_ _07783_ vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__a221o_1
X_14890_ net1090 _08419_ vssd1 vssd1 vccd1 vccd1 _08667_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout64_X net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17270__A1 _02275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10893__A1 game.CPU.applesa.ab.XMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ game.writer.tracker.frame\[522\] net842 net834 game.writer.tracker.frame\[521\]
+ vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__o22a_1
XFILLER_0_202_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_241_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11942__X _05830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16560_ net1889 _02481_ _02487_ net125 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[83\]
+ sky130_fd_sc_hd__a22o_1
X_13772_ game.writer.tracker.frame\[158\] net844 net838 game.writer.tracker.frame\[157\]
+ vssd1 vssd1 vccd1 vccd1 _07646_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10984_ _04862_ _04863_ _04864_ _04868_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__or4_1
XANTENNA__16229__Y _02237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15511_ net888 _01532_ _01531_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_167_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12723_ game.writer.tracker.frame\[100\] game.writer.tracker.frame\[101\] net995
+ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16491_ net199 _02315_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_256_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09779__B net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13081__S net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09131__Y _03380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18230_ net649 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__inv_2
X_15442_ _01468_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ _06246_ _06452_ _06529_ _06530_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__nand4_2
XFILLER_0_242_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_178_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11605_ net745 _05490_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18161_ net631 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__inv_2
XANTENNA__15797__A game.CPU.applesa.ab.absxs.body_y\[50\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15373_ _08878_ _08883_ game.writer.updater.commands.cmd_num\[0\] vssd1 vssd1 vccd1
+ vccd1 _08915_ sky130_fd_sc_hd__mux2_1
X_12585_ game.CPU.applesa.ab.absxs.body_y\[8\] net361 vssd1 vssd1 vccd1 vccd1 _06462_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__17325__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17112_ _02359_ _02693_ net734 vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__o21a_1
X_11536_ net790 net249 vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_133_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14324_ game.CPU.applesa.ab.absxs.body_x\[75\] net1046 vssd1 vssd1 vccd1 vccd1 _08198_
+ sky130_fd_sc_hd__or2_1
X_18092_ net591 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__inv_2
XANTENNA__11070__B2 game.CPU.applesa.ab.absxs.body_y\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11740__A1_N _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_312_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13347__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17043_ _02398_ net85 _02684_ net1656 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[369\]
+ sky130_fd_sc_hd__a22o_1
X_14255_ _08122_ _08124_ _08125_ _08128_ vssd1 vssd1 vccd1 vccd1 _08129_ sky130_fd_sc_hd__or4_2
XFILLER_0_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11467_ net565 _05351_ _05350_ net744 vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_150_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13898__A1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ net496 _07079_ net684 vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13898__B2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17089__B2 game.writer.tracker.frame\[401\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10418_ game.CPU.down_button.eD1.Q2 game.CPU.down_button.eD1.Q1 vssd1 vssd1 vccd1
+ vccd1 _04563_ sky130_fd_sc_hd__nand2b_2
X_14186_ _03284_ net1072 net873 game.CPU.applesa.ab.absxs.body_x\[19\] vssd1 vssd1
+ vccd1 vccd1 _08060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11398_ net567 _05282_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_267_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16836__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11373__A2 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13137_ game.writer.tracker.frame\[162\] game.writer.tracker.frame\[163\] net1005
+ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_209_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ game.CPU.walls.rand_wall.counter2\[3\] game.CPU.walls.rand_wall.counter2\[2\]
+ game.CPU.walls.rand_wall.counter2\[1\] game.CPU.walls.rand_wall.counter2\[0\] vssd1
+ vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_280_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18994_ net1197 _00220_ _00665_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[39\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_264_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13068_ _06938_ _06939_ _06941_ _06940_ net491 net686 vssd1 vssd1 vccd1 vccd1 _06942_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10381__A1_N net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17945_ net651 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__inv_2
XFILLER_0_209_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11565__A game.CPU.applesa.ab.check_walls.above.walls\[135\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ game.CPU.applesa.ab.check_walls.above.walls\[45\] net388 vssd1 vssd1 vccd1
+ vccd1 _05906_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_224_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17876_ net636 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__inv_2
X_19615_ clknet_leaf_21_clk game.writer.tracker.next_frame\[210\] net1336 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[210\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_283_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17261__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09035__A game.CPU.applesa.ab.absxs.body_x\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16827_ net156 _02365_ net98 net715 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__o31a_1
XFILLER_0_250_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_348_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19546_ clknet_leaf_49_clk game.writer.tracker.next_frame\[141\] net1297 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[141\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16758_ game.writer.tracker.frame\[180\] _02588_ vssd1 vssd1 vccd1 vccd1 _02589_
+ sky130_fd_sc_hd__and2_1
XANTENNA__13822__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_278_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15709_ game.CPU.applesa.ab.absxs.body_y\[8\] net452 vssd1 vssd1 vccd1 vccd1 _01721_
+ sky130_fd_sc_hd__xnor2_1
X_19477_ clknet_leaf_20_clk game.writer.tracker.next_frame\[72\] net1315 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[72\] sky130_fd_sc_hd__dfrtp_1
X_16689_ _02464_ net62 _02563_ net1951 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[136\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18917__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_291_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09230_ game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1 vssd1 vccd1 vccd1
+ _03479_ sky130_fd_sc_hd__inv_2
X_18428_ net586 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__inv_2
XFILLER_0_347_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14378__A2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_233_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__B game.CPU.applesa.ab.absxs.body_x\[54\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_118_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_319_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09161_ game.CPU.applesa.ab.check_walls.above.walls\[56\] vssd1 vssd1 vccd1 vccd1
+ _03410_ sky130_fd_sc_hd__inv_2
X_18359_ net597 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18083__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16155__X _02167_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15500__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_303_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09092_ game.CPU.applesa.ab.absxs.body_y\[49\] vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload50_A clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16524__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13939__B game.CPU.applesa.ab.check_walls.above.walls\[65\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11299__X _05189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_302_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_330_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout111_A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10644__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13433__S0 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14116__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_309_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout209_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_275_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16827__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13955__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1020_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09994_ game.CPU.apple_location\[5\] net1494 _04207_ vssd1 vssd1 vccd1 vccd1 _01370_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_244_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ net1105 vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout480_A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16050__B net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_327_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13510__B1 _07383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout199_X net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__A game.CPU.applesa.ab.check_walls.above.walls\[51\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17252__A1 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_230_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18258__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout745_A _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17004__A1 _02328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18597__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11922__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_338_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout912_A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19842__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1275_X net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16212__C1 _01814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09428_ net1082 _03441_ _03442_ net1135 vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_338_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15113__C game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09359_ net1108 game.CPU.applesa.ab.check_walls.above.walls\[192\] vssd1 vssd1 vccd1
+ vccd1 _03602_ sky130_fd_sc_hd__xor2_1
XANTENNA__16506__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13672__S0 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_306_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12370_ game.CPU.applesa.ab.absxs.body_x\[115\] net530 vssd1 vssd1 vccd1 vccd1 _06247_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__16515__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19992__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_288_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_185_Right_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11321_ net563 _04775_ _05209_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__o21a_2
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ net1053 _03440_ _03443_ net938 vssd1 vssd1 vccd1 vccd1 _07914_ sky130_fd_sc_hd__o22a_1
X_11252_ game.CPU.applesa.ab.absxs.body_x\[115\] net545 net409 game.CPU.applesa.ab.absxs.body_x\[114\]
+ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_344_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19222__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ _04395_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11183_ game.CPU.applesa.ab.absxs.body_x\[84\] net326 vssd1 vssd1 vccd1 vccd1 _05073_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__16294__A2 _08400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17491__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ game.CPU.randy.f1.c1.count\[5\] game.CPU.randy.f1.c1.count\[7\] _04327_ _04328_
+ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__or4_1
XFILLER_0_207_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15991_ game.CPU.applesa.ab.check_walls.above.walls\[103\] net432 vssd1 vssd1 vccd1
+ vccd1 _02003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_261_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17730_ game.CPU.applesa.ab.count_luck\[6\] game.CPU.applesa.ab.count_luck\[5\] _03093_
+ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__and3_1
X_10065_ net1144 _04218_ _04221_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__o21ba_1
X_14942_ _08676_ _08683_ _08718_ vssd1 vssd1 vccd1 vccd1 _08719_ sky130_fd_sc_hd__nor3_1
XANTENNA__19372__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17243__B2 game.writer.tracker.frame\[512\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17661_ game.CPU.kyle.L1.cnt_500hz\[9\] game.CPU.kyle.L1.cnt_500hz\[10\] game.CPU.kyle.L1.cnt_500hz\[11\]
+ _03047_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__and4_1
XFILLER_0_89_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14873_ game.CPU.walls.abc.number\[5\] game.CPU.walls.abc.number\[1\] game.CPU.walls.abc.counter
+ vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_242_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19400_ clknet_leaf_47_clk _01400_ net1298 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.x\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_106_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16612_ net2004 _02515_ _02521_ _02522_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[100\]
+ sky130_fd_sc_hd__a22o_1
X_13824_ _07668_ _07681_ _07697_ net177 vssd1 vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17592_ game.CPU.kyle.L1.cnt_20ms\[1\] game.CPU.kyle.L1.cnt_20ms\[0\] game.CPU.kyle.L1.cnt_20ms\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19331_ clknet_leaf_72_clk net1431 _00936_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twomode.number\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_159_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16543_ net1723 _02474_ _02475_ net124 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[78\]
+ sky130_fd_sc_hd__a22o_1
X_13755_ game.writer.tracker.frame\[161\] game.writer.tracker.frame\[163\] game.writer.tracker.frame\[164\]
+ game.writer.tracker.frame\[162\] net969 net1005 vssd1 vssd1 vccd1 vccd1 _07629_
+ sky130_fd_sc_hd__mux4_1
X_10967_ net1265 net406 vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__or2_1
XFILLER_0_174_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ _06554_ _06564_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__nor2_1
X_19262_ clknet_leaf_9_clk _00050_ _00892_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_329_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16474_ net167 _02342_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__nand2_8
XANTENNA__15023__C game.CPU.applesa.ab.check_walls.above.walls\[51\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13686_ game.writer.tracker.frame\[481\] game.writer.tracker.frame\[483\] game.writer.tracker.frame\[484\]
+ game.writer.tracker.frame\[482\] net974 net1010 vssd1 vssd1 vccd1 vccd1 _07560_
+ sky130_fd_sc_hd__mux4_1
X_10898_ game.CPU.applesa.ab.check_walls.collision_down _04798_ _04799_ vssd1 vssd1
+ vccd1 vccd1 _04800_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_344_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13568__A0 game.writer.tracker.frame\[329\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18213_ net666 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
X_15425_ _01438_ _01451_ _01452_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__a21bo_1
X_19193_ clknet_leaf_54_clk net341 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.y_final\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12637_ _06398_ _06400_ _06401_ _06513_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18144_ net631 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__inv_2
XFILLER_0_288_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15356_ _08883_ _08897_ vssd1 vssd1 vccd1 vccd1 _08898_ sky130_fd_sc_hd__and2_1
X_12568_ game.CPU.applesa.ab.absxs.body_y\[117\] net524 vssd1 vssd1 vccd1 vccd1 _06445_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_331_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_215_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14307_ _03247_ net1045 net959 _03315_ _08176_ vssd1 vssd1 vccd1 vccd1 _08181_ sky130_fd_sc_hd__a221o_1
X_11519_ net831 net262 _05395_ _05406_ _05407_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18075_ net657 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__inv_2
X_12499_ game.CPU.applesa.ab.absxs.body_y\[61\] net525 vssd1 vssd1 vccd1 vccd1 _06376_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__12008__X _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15287_ _08815_ _08837_ _08838_ _08812_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a22o_1
Xhold207 game.writer.tracker.frame\[493\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xwire193 _05405_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_1
Xhold218 game.writer.tracker.frame\[342\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 game.writer.tracker.frame\[371\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ _02365_ _02670_ net717 vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__o21a_1
XFILLER_0_300_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14238_ game.CPU.applesa.ab.absxs.body_x\[114\] net1056 vssd1 vssd1 vccd1 vccd1 _08112_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__15974__B net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_296_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ game.CPU.applesa.ab.absxs.body_y\[105\] net964 vssd1 vssd1 vccd1 vccd1 _08043_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_298_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout709 _06594_ vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19715__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18977_ net1196 _00202_ _00648_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10911__B _04808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_265_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17928_ net606 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__inv_2
XFILLER_0_294_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1280 net1281 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__clkbuf_4
Xfanout1291 net1292 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_280_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17859_ game.writer.updater.commands.count\[12\] _03178_ _03181_ _03175_ vssd1 vssd1
+ vccd1 vccd1 _01421_ sky130_fd_sc_hd__o211a_1
XFILLER_0_212_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_201_Left_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19865__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11582__X _05471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19529_ clknet_leaf_22_clk game.writer.tracker.next_frame\[124\] net1344 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[124\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_287_Right_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10609__B2 game.CPU.applesa.ab.absxs.body_x\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09475__A1 net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09475__B2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_313_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_307_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13559__B1 net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09213_ game.CPU.applesa.ab.check_walls.above.walls\[158\] vssd1 vssd1 vccd1 vccd1
+ _03462_ sky130_fd_sc_hd__inv_2
XFILLER_0_335_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_315_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13654__S0 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout326_A game.CPU.applesa.ab.absxs.next_head\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16760__A3 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1068_A game.CPU.applesa.x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1 vccd1 vccd1
+ _03393_ sky130_fd_sc_hd__inv_2
XANTENNA__13669__B _07488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09075_ game.CPU.applesa.ab.absxs.body_y\[108\] vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__inv_2
XANTENNA__10374__A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout114_X net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18541__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16512__A3 _02454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1235_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14523__A2 _07742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15884__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout695_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13731__B1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_338_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout862_A net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ net1158 net1262 vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_283_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_164_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16028__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18984__Q game.CPU.applesa.ab.check_walls.above.walls\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13624__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11933__A game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11870_ net831 net312 net393 net832 _05757_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__o221a_1
XFILLER_0_354_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13798__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10821_ game.CPU.applesa.ab.absxs.body_y\[8\] _04689_ _04707_ game.CPU.applesa.ab.absxs.body_y\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_254_Right_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17528__A2 _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09897__X _04140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13540_ game.writer.tracker.frame\[119\] net710 net673 game.writer.tracker.frame\[120\]
+ _07413_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__o221a_1
X_10752_ game.CPU.applesa.ab.absxs.body_y\[111\] _04665_ _04666_ game.CPU.applesa.ab.absxs.body_y\[107\]
+ vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_253_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12470__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_326_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10268__B net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16200__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13471_ _07343_ _07344_ net214 vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_175_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10683_ game.CPU.applesa.ab.absxs.body_x\[9\] _04689_ _04707_ game.CPU.applesa.ab.absxs.body_x\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__a22o_1
XFILLER_0_353_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16236__A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_350_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_299_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15210_ _08777_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__inv_2
XANTENNA__15140__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ game.CPU.applesa.ab.absxs.body_x\[33\] net375 net517 game.CPU.applesa.ab.absxs.body_y\[34\]
+ _06297_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__a221o_1
X_16190_ _01635_ _02125_ _02127_ _02128_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_117_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15141_ net1209 net1235 game.CPU.applesa.ab.check_walls.above.walls\[169\] vssd1
+ vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__and3_1
X_12353_ game.CPU.applesa.ab.absxs.body_y\[79\] net367 vssd1 vssd1 vccd1 vccd1 _06230_
+ sky130_fd_sc_hd__or2_1
X_11304_ game.CPU.applesa.ab.apple_possible\[6\] _05192_ vssd1 vssd1 vccd1 vccd1 _05193_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_132_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19738__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15072_ net1212 net1238 game.CPU.applesa.ab.check_walls.above.walls\[100\] vssd1
+ vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__and3_1
XFILLER_0_294_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11099__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14514__A2 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12284_ game.CPU.applesa.ab.check_walls.above.walls\[134\] net417 vssd1 vssd1 vccd1
+ vccd1 _06170_ sky130_fd_sc_hd__xnor2_1
XANTENNA__20045__X net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14023_ net856 net786 game.CPU.applesa.ab.check_walls.above.walls\[161\] net881 vssd1
+ vssd1 vccd1 vccd1 _07897_ sky130_fd_sc_hd__a2bb2o_1
X_18900_ clknet_leaf_68_clk _01267_ _00584_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.good_collision
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13722__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17067__A _02240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11235_ game.CPU.applesa.ab.absxs.body_x\[12\] net415 vssd1 vssd1 vccd1 vccd1 _05125_
+ sky130_fd_sc_hd__xnor2_1
X_19880_ clknet_leaf_25_clk game.writer.tracker.next_frame\[475\] net1319 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[475\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10571__X _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_264_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10536__B1 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_293_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_248_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16402__C net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18831_ clknet_leaf_0_clk _01222_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11166_ _05053_ _05054_ _05055_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_112_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19888__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18762__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10117_ _04318_ game.CPU.applesa.apple_location2_n\[2\] _04311_ vssd1 vssd1 vccd1
+ vccd1 _01342_ sky130_fd_sc_hd__mux2_1
X_18762_ clknet_leaf_50_clk _01179_ _00499_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[60\]
+ sky130_fd_sc_hd__dfrtp_4
X_11097_ _03270_ net406 vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__xnor2_1
X_15974_ game.CPU.applesa.ab.absxs.body_x\[67\] net463 vssd1 vssd1 vccd1 vccd1 _01986_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_128_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_303_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17216__A1 _02238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17713_ game.CPU.applesa.ab.count_luck\[0\] _03084_ vssd1 vssd1 vccd1 vccd1 _03086_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_262_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10048_ net1271 net846 vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__nor2_4
X_14925_ _08678_ _08681_ _08682_ _08679_ vssd1 vssd1 vccd1 vccd1 _08702_ sky130_fd_sc_hd__o31a_1
XFILLER_0_264_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18693_ clknet_leaf_58_clk _01110_ _00430_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[35\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_215_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold90 game.CPU.applesa.apple_location2_n\[3\] vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
X_17644_ game.CPU.kyle.L1.cnt_500hz\[3\] game.CPU.kyle.L1.cnt_500hz\[4\] _08801_ game.CPU.kyle.L1.cnt_500hz\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__a31o_1
XFILLER_0_264_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14856_ _08647_ _08648_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[11\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09313__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13807_ net279 _07674_ _07680_ net247 vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_201_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09457__A1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17575_ _02858_ _02964_ _02994_ _02998_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_221_Right_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14787_ _03512_ _08603_ vssd1 vssd1 vccd1 vccd1 _08606_ sky130_fd_sc_hd__nor2_1
XANTENNA__09457__B2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_275_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ _05874_ _05875_ _05876_ _05885_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__o31a_1
XFILLER_0_280_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19314_ net1164 _00038_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.out_random_2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16526_ _02286_ net144 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__nor2_2
XFILLER_0_187_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11264__A1 game.CPU.applesa.ab.absxs.body_y\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13738_ game.writer.tracker.frame\[209\] game.writer.tracker.frame\[211\] game.writer.tracker.frame\[212\]
+ game.writer.tracker.frame\[210\] net978 net1026 vssd1 vssd1 vccd1 vccd1 _07612_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_217_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15969__B net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_280_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19245_ clknet_leaf_17_clk _00059_ _00883_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__19268__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16457_ _02234_ _02277_ _02413_ net733 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__o31a_1
X_13669_ net183 _07488_ _07504_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__and3_1
XANTENNA__14218__X _08092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_344_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13122__X _06996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15050__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15408_ game.writer.updater.commands.cmd_num\[2\] game.writer.updater.commands.cmd_num\[3\]
+ game.writer.updater.commands.cmd_num\[4\] vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__or3b_2
X_19176_ clknet_leaf_4_clk _01295_ _00838_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_16388_ _02362_ net165 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__and2b_4
XFILLER_0_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15985__A game.CPU.applesa.ab.check_walls.above.walls\[70\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_18127_ net578 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__inv_2
XANTENNA__13961__B1 game.CPU.applesa.ab.check_walls.above.walls\[179\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_332_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15339_ game.writer.updater.commands.cmd_num\[1\] game.writer.updater.commands.cmd_num\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08881_ sky130_fd_sc_hd__nand2_1
XANTENNA__10194__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14505__A2 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18058_ net632 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_285_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_257_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11319__A2 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17009_ _02498_ net84 _02674_ net1805 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[345\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_257_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09900_ _03755_ _03758_ _03763_ _03868_ _04142_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__o311a_1
XANTENNA__10790__A3 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_286_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10922__A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__B1 _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16258__A2 _06573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_228_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17455__A1 _03197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20020_ net1276 vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
X_09831_ _04069_ _04070_ _04073_ _04068_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__a211o_1
Xfanout517 _06214_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_4
Xfanout528 net532 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__buf_4
XFILLER_0_284_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14269__A1 game.CPU.applesa.ab.absxs.body_x\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkload13_A clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout539 net540 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_356_Right_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14269__B2 game.CPU.applesa.ab.absxs.body_y\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09762_ _04000_ _04001_ _04002_ _04004_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__a211o_1
X_09693_ net1084 game.CPU.applesa.ab.absxs.body_x\[7\] vssd1 vssd1 vccd1 vccd1 _03936_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__09696__A1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09696__B2 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13444__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout276_A _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_339_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_317_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12568__B net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09223__A game.CPU.applesa.ab.check_walls.above.walls\[171\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09448__A1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09448__B2 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout443_A _08429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16981__A3 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_239_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15879__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout610_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1352_A net1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout708_A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18635__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_340_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_323_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09127_ net943 vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1140_X net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18271__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09620__B2 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1238_X net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16497__A2 _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09058_ game.CPU.applesa.ab.absxs.body_y\[53\] vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__inv_2
XANTENNA__18979__Q game.CPU.applesa.ab.check_walls.above.walls\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_328_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_276_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13704__A0 game.writer.tracker.frame\[497\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_107_Left_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18785__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 game.writer.tracker.frame\[82\] vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17318__C _02413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 game.writer.tracker.frame\[539\] vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 game.writer.tracker.frame\[85\] vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ game.CPU.applesa.ab.absxs.body_y\[89\] net543 vssd1 vssd1 vccd1 vccd1 _04910_
+ sky130_fd_sc_hd__xnor2_1
Xhold593 game.CPU.applesa.apple_location2_n\[0\] vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11191__B1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_323_Right_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_216_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12971_ net509 _06844_ _06843_ net211 vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__o211a_1
XANTENNA__09687__A1 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13354__S net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_271_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15135__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14710_ net55 _08546_ _08547_ vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__and3_1
X_11922_ net781 net311 vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__xor2_1
X_15690_ game.CPU.applesa.ab.absxs.body_y\[7\] net433 vssd1 vssd1 vccd1 vccd1 _01702_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_339_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_Left_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14641_ game.CPU.clock1.counter\[18\] game.CPU.clock1.counter\[19\] _08479_ game.CPU.clock1.counter\[20\]
+ vssd1 vssd1 vccd1 vccd1 _08483_ sky130_fd_sc_hd__a31o_1
X_11853_ _03435_ net312 vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19410__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18446__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14432__B2 game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_345_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17360_ net1116 _08748_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__or2_1
X_10804_ game.CPU.applesa.ab.absxs.body_y\[25\] _04695_ _04698_ game.CPU.applesa.ab.absxs.body_y\[21\]
+ vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__a22o_1
XANTENNA__16709__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12443__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14572_ net1264 _08432_ _08434_ _00039_ vssd1 vssd1 vccd1 vccd1 game.CPU.state1.Qn\[1\]
+ sky130_fd_sc_hd__a22o_1
X_11784_ game.CPU.applesa.ab.check_walls.above.walls\[39\] net312 vssd1 vssd1 vccd1
+ vccd1 _05672_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11246__B2 game.CPU.applesa.ab.absxs.body_y\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15789__B net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_345_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16311_ net236 _02307_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__nand2_2
XFILLER_0_82_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_306_Left_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13523_ net186 _07391_ _07396_ net177 vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__o211a_1
XFILLER_0_184_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17291_ net175 net116 _02364_ _02753_ net1498 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[547\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_103_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10735_ game.CPU.applesa.ab.absxs.body_y\[20\] _04645_ _04652_ game.CPU.applesa.ab.absxs.body_y\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13618__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16185__B2 game.CPU.applesa.ab.check_walls.above.walls\[106\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19030_ net1193 _00260_ _00701_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[75\]
+ sky130_fd_sc_hd__dfrtp_4
X_16242_ net274 _02226_ _02227_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14196__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19560__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13454_ net689 _07027_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__or2_1
XFILLER_0_250_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10666_ game.CPU.applesa.ab.absxs.body_x\[19\] _04699_ _04700_ game.CPU.applesa.ab.absxs.body_x\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__a22o_1
XFILLER_0_353_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12746__A1 game.writer.tracker.frame\[81\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ game.CPU.applesa.ab.absxs.body_x\[54\] net373 vssd1 vssd1 vccd1 vccd1 _06282_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13385_ _06862_ _06883_ net679 vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__mux2_1
X_16173_ _03276_ net353 game.CPU.walls.rand_wall.abduyd.next_wall\[7\] _03345_ _02184_
+ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a221o_1
XANTENNA__17134__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09611__A1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10597_ _03230_ net263 vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__nor2_1
XANTENNA__09611__B2 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Left_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15124_ net1208 net1233 game.CPU.applesa.ab.check_walls.above.walls\[152\] vssd1
+ vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17068__Y _02692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12336_ _04226_ _04258_ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_267_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19932_ clknet_leaf_48_clk game.writer.tracker.next_frame\[527\] net1302 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[527\] sky130_fd_sc_hd__dfrtp_1
X_12267_ _05930_ _05931_ _06151_ _06152_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__and4b_1
X_15055_ net1217 net1245 game.CPU.applesa.ab.check_walls.above.walls\[83\] vssd1 vssd1
+ vccd1 vccd1 _00278_ sky130_fd_sc_hd__and3_1
XANTENNA__10509__B1 _04626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10742__A game.CPU.applesa.ab.absxs.body_y\[106\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13171__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14006_ net877 game.CPU.applesa.ab.check_walls.above.walls\[138\] _03453_ net1043
+ vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__a22o_1
X_11218_ _03246_ net324 vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_315_Left_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19863_ clknet_leaf_20_clk game.writer.tracker.next_frame\[458\] net1315 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[458\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09308__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12198_ game.CPU.applesa.ab.check_walls.above.walls\[53\] net549 vssd1 vssd1 vccd1
+ vccd1 _06084_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15029__B net1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11721__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18814_ clknet_leaf_72_clk game.CPU.clock1.next_counter\[17\] _00551_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[17\] sky130_fd_sc_hd__dfrtp_1
X_11149_ _03260_ net546 vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__nand2_1
X_19794_ clknet_leaf_36_clk game.writer.tracker.next_frame\[389\] net1355 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[389\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13459__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16660__A2 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18745_ clknet_leaf_10_clk _01162_ _00482_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_222_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15957_ game.CPU.applesa.ab.check_walls.above.walls\[24\] net356 vssd1 vssd1 vccd1
+ vccd1 _01969_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09678__A1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Left_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09678__B2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_223_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14908_ net1171 _08426_ _08424_ game.CPU.applesa.ab.YMAX\[0\] vssd1 vssd1 vccd1 vccd1
+ _08685_ sky130_fd_sc_hd__o211a_1
XFILLER_0_163_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18676_ clknet_leaf_8_clk _01093_ _00413_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16948__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15888_ game.CPU.applesa.ab.check_walls.above.walls\[136\] net354 vssd1 vssd1 vccd1
+ vccd1 _01900_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12388__B game.CPU.applesa.twoapples.absxs.next_head\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09043__A game.CPU.applesa.ab.absxs.body_x\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17627_ game.CPU.kyle.L1.cnt_20ms\[15\] _03032_ net577 vssd1 vssd1 vccd1 vccd1 _03033_
+ sky130_fd_sc_hd__a21oi_1
X_14839_ game.CPU.randy.f1.c1.count\[5\] game.CPU.randy.f1.c1.count\[4\] _08635_ vssd1
+ vssd1 vccd1 vccd1 _08638_ sky130_fd_sc_hd__and3_1
XANTENNA__10189__A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14884__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13857__S0 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_330_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_76 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_324_Left_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09978__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18658__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17558_ _02849_ _02923_ _02965_ _02850_ _02858_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12434__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19903__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16509_ net150 net128 _02452_ _02446_ net1530 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[67\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_156_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17489_ _02781_ _02784_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10917__A net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19228_ clknet_leaf_57_clk net1422 _00866_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.normal1.number\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14187__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_312_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_288_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13934__B1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19159_ clknet_leaf_3_clk _01280_ _00830_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.counter2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17125__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16163__X _02175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16604__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_258_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17140__A3 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16323__B net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13439__S net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_333_Left_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_285_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14124__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17428__A1 net1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout303 net304 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_4
Xfanout314 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_4
Xfanout325 net326 vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16610__Y _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20003_ clknet_leaf_44_clk game.writer.updater.update.next\[1\] net1300 vssd1 vssd1
+ vccd1 vccd1 game.writer.updater.commands.mode\[1\] sky130_fd_sc_hd__dfrtp_2
Xfanout336 net340 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_6
X_09814_ net1098 _03280_ game.CPU.applesa.ab.absxs.body_y\[26\] net903 vssd1 vssd1
+ vccd1 vccd1 _04057_ sky130_fd_sc_hd__a22o_1
Xfanout347 game.CPU.walls.rand_wall.abduyd.next_wall\[2\] vssd1 vssd1 vccd1 vccd1
+ net347 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_323_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout369 game.CPU.applesa.twoapples.absxs.next_head\[5\] vssd1 vssd1 vccd1 vccd1
+ net369 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1100_A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16651__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ net1087 _03417_ net815 net899 _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__a221o_1
XANTENNA__19433__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12579__A game.CPU.applesa.ab.absxs.body_x\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_335_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16939__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ net909 game.CPU.applesa.ab.absxs.body_y\[103\] vssd1 vssd1 vccd1 vccd1 _03919_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12298__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16338__X _02328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1090_X net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18266__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout825_A game.CPU.applesa.ab.check_walls.above.walls\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14414__A1 game.CPU.applesa.ab.absxs.body_x\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_221_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1188_X net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14414__B2 game.CPU.applesa.ab.absxs.body_x\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_327_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_355_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19583__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14965__A2 game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19540__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16167__A1 game.CPU.applesa.ab.absxs.body_y\[76\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10520_ net933 game.CPU.applesa.ab.absxs.body_x\[58\] vssd1 vssd1 vccd1 vccd1 _04634_
+ sky130_fd_sc_hd__and2_1
XANTENNA__16217__C net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15121__C game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10451_ _04579_ _04585_ _04578_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_323_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13170_ net231 _07039_ net280 vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__a21o_1
X_10382_ net1125 _03203_ game.CPU.apple_location2\[2\] net919 _04528_ vssd1 vssd1
+ vccd1 vccd1 _04535_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout982_X net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_288_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12121_ game.CPU.applesa.ab.check_walls.above.walls\[173\] net387 vssd1 vssd1 vccd1
+ vccd1 _06008_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13689__C1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14034__A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09128__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14350__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ _05936_ _05937_ _05938_ _05935_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__a211o_1
Xhold390 game.writer.tracker.frame\[499\] vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_261_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11003_ _04887_ _04888_ _04891_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__or4_1
XANTENNA__13873__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16860_ net133 _02412_ net122 _02625_ net1521 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[245\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_183_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08967__A game.CPU.applesa.ab.absxs.body_y\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 net871 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_4
X_15811_ _01817_ _01818_ _01820_ _01821_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__or4_1
Xfanout881 net882 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_8
X_16791_ _02470_ net102 _02598_ net1605 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[203\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_217_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout892 net896 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_125_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18530_ net601 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__inv_2
X_15742_ game.CPU.applesa.ab.check_walls.above.walls\[175\] net430 vssd1 vssd1 vccd1
+ vccd1 _01754_ sky130_fd_sc_hd__nor2_1
X_12954_ _06757_ _06760_ net680 vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__mux2_1
XANTENNA__12664__B1 _06540_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__B2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13861__C1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18800__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19628__RESET_B net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19926__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18461_ net652 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__inv_2
X_11905_ net805 net302 _05792_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__a21bo_1
X_15673_ game.CPU.applesa.ab.check_walls.above.walls\[10\] net348 vssd1 vssd1 vccd1
+ vccd1 _01685_ sky130_fd_sc_hd__or2_1
XFILLER_0_319_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12885_ game.writer.tracker.frame\[10\] game.writer.tracker.frame\[11\] net1002 vssd1
+ vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__mux2_1
XANTENNA__12001__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17412_ _02839_ _02841_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__nand2_1
XFILLER_0_212_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14624_ net2009 _08470_ _08472_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[13\]
+ sky130_fd_sc_hd__a21oi_1
X_11836_ game.CPU.applesa.ab.check_walls.above.walls\[149\] net305 vssd1 vssd1 vccd1
+ vccd1 _05724_ sky130_fd_sc_hd__xor2_1
X_18392_ net600 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_346_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_272_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12967__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16408__B _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17343_ game.CPU.kyle.L1.nextState\[5\] game.CPU.kyle.L1.nextState\[4\] game.CPU.kyle.L1.nextState\[2\]
+ game.CPU.kyle.L1.nextState\[3\] vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__or4b_4
XFILLER_0_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14555_ net458 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.abduyd.next_wall\[3\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__18950__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ _05645_ _05647_ _05654_ _05644_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_194_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ net278 _07312_ _07320_ net241 vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__a211o_2
XFILLER_0_125_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17274_ net176 _02258_ net69 _02749_ net1802 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[535\]
+ sky130_fd_sc_hd__a32o_1
X_10718_ game.CPU.applesa.ab.absxs.body_y\[52\] _04609_ _04637_ game.CPU.applesa.ab.absxs.body_y\[48\]
+ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14486_ _08213_ _08220_ _08345_ _08184_ _08117_ vssd1 vssd1 vccd1 vccd1 _08360_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11698_ game.CPU.applesa.ab.check_walls.above.walls\[162\] net766 vssd1 vssd1 vccd1
+ vccd1 _05587_ sky130_fd_sc_hd__xor2_2
XFILLER_0_36_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19013_ net1196 _00241_ _00684_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[58\]
+ sky130_fd_sc_hd__dfrtp_4
X_16225_ net175 _02231_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__nor2_2
X_13437_ _06939_ _06941_ _06956_ _06940_ net702 net491 vssd1 vssd1 vccd1 vccd1 _07311_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_341_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10649_ _04693_ game.CPU.applesa.ab.absxs.body_x\[41\] _04690_ vssd1 vssd1 vccd1
+ vccd1 _01112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19306__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16156_ _01646_ _01648_ _01650_ _01651_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__or4_1
X_13368_ _06679_ _06681_ _06690_ _06680_ net693 net478 vssd1 vssd1 vccd1 vccd1 _07242_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17122__A3 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15107_ net1203 net1229 game.CPU.applesa.ab.check_walls.above.walls\[135\] vssd1
+ vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__and3_1
XANTENNA__10745__A3 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ _06108_ _06111_ _06173_ _06180_ _06192_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__o2111a_1
X_16087_ game.CPU.applesa.ab.check_walls.above.walls\[147\] net459 net439 game.CPU.applesa.ab.check_walls.above.walls\[150\]
+ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a2bb2o_1
X_13299_ _06752_ _06780_ _06781_ _06782_ net513 net706 vssd1 vssd1 vccd1 vccd1 _07173_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_294_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_283_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_35_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19915_ clknet_leaf_24_clk game.writer.tracker.next_frame\[510\] net1339 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[510\] sky130_fd_sc_hd__dfrtp_1
X_15038_ net1221 net1247 game.CPU.applesa.ab.check_walls.above.walls\[66\] vssd1 vssd1
+ vccd1 vccd1 _00259_ sky130_fd_sc_hd__and3_1
XANTENNA__14341__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_225_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19456__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_280_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_299_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19846_ clknet_leaf_40_clk game.writer.tracker.next_frame\[441\] net1357 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[441\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10902__B1 _04796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_142_Left_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16633__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19777_ clknet_leaf_26_clk game.writer.tracker.next_frame\[372\] net1312 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[372\] sky130_fd_sc_hd__dfrtp_1
X_16989_ _02471_ net88 _02667_ net1554 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[332\]
+ sky130_fd_sc_hd__a22o_1
X_09530_ _03770_ _03771_ _03772_ _03766_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__a211o_1
X_18728_ clknet_leaf_13_clk _01145_ _00465_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[110\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13852__C1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _03698_ _03699_ _03703_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__or3b_2
X_18659_ clknet_leaf_59_clk _01076_ _00396_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[77\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16397__B2 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16158__X _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18086__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_305_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15503__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_294_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12407__B1 game.CPU.applesa.twoapples.absxs.next_head\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09392_ net914 game.CPU.applesa.ab.check_walls.above.walls\[161\] game.CPU.applesa.ab.check_walls.above.walls\[163\]
+ net925 _03632_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__a221o_1
XFILLER_0_337_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12958__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_236_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09501__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11750__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16149__A1 _01725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_151_Left_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout239_A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13958__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1050_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_A net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_341_Left_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13383__A1 _07209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1148_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_258_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12581__B net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_325_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11478__A game.CPU.applesa.ab.check_walls.above.walls\[49\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1315_A net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11197__B net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16872__A2 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_247_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15892__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout100 _02559_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__buf_4
Xfanout111 net112 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout775_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 net1113 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_4
Xfanout122 _02597_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_4
XFILLER_0_245_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout133 _02235_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_4
Xfanout144 _02440_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12894__A0 game.writer.tracker.frame\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1103_X net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout155 _02270_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_2
Xfanout166 _02363_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_4
XANTENNA__16085__B1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18823__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_346_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19949__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout177 _06639_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout188 net189 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_4
Xfanout199 _02288_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_2
XANTENNA_fanout942_A game.CPU.applesa.y\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14301__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19792__RESET_B net1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ net1107 game.CPU.applesa.ab.absxs.body_x\[32\] vssd1 vssd1 vccd1 vccd1 _03971_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_241_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_241_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_336_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _03894_ _03895_ _03900_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__a211o_1
XANTENNA__18973__CLK net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11845__A2_N net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12670_ game.writer.updater.commands.mode\[1\] game.writer.updater.commands.mode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16228__B net141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09411__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15132__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11621_ game.CPU.applesa.ab.check_walls.above.walls\[185\] net770 vssd1 vssd1 vccd1
+ vccd1 _05510_ sky130_fd_sc_hd__xor2_1
XFILLER_0_194_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_239_Left_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09814__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10557__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09814__B2 net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19329__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14340_ game.CPU.applesa.ab.absxs.body_y\[38\] net951 vssd1 vssd1 vccd1 vccd1 _08214_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_231_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11552_ game.CPU.applesa.ab.check_walls.above.walls\[194\] net767 vssd1 vssd1 vccd1
+ vccd1 _05441_ sky130_fd_sc_hd__xor2_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10503_ game.CPU.applesa.ab.absxs.body_x\[78\] _04623_ _04624_ game.CPU.applesa.ab.absxs.body_x\[74\]
+ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__a22o_1
X_14271_ _03341_ net962 net858 game.CPU.applesa.ab.absxs.body_y\[51\] _08144_ vssd1
+ vssd1 vccd1 vccd1 _08145_ sky130_fd_sc_hd__o221a_1
X_11483_ net567 _05366_ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16560__B2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16244__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_311_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16010_ game.CPU.applesa.ab.absxs.body_y\[61\] net446 vssd1 vssd1 vccd1 vccd1 _02022_
+ sky130_fd_sc_hd__xnor2_1
X_13222_ game.writer.tracker.frame\[392\] game.writer.tracker.frame\[393\] net1036
+ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__mux2_1
X_10434_ game.CPU.applesa.ab.absxs.body_x\[7\] net847 _04158_ net1449 vssd1 vssd1
+ vccd1 vccd1 _01210_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_347_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12491__B net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19479__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13079__S net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_249_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11924__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13153_ game.writer.tracker.frame\[178\] game.writer.tracker.frame\[179\] net1035
+ vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10365_ net2020 _04526_ _04525_ _04518_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13126__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ net796 net295 net292 net797 vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__o2bb2a_1
X_13084_ net477 _06957_ net683 vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__a21o_1
X_17961_ net657 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__inv_2
X_10296_ net851 game.CPU.applesa.ab.good_spot_next game.CPU.applesa.ab.apple_location\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16250__Y _02258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13677__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16912_ _02327_ net95 _02646_ net1798 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[276\]
+ sky130_fd_sc_hd__a22o_1
X_19700_ clknet_leaf_30_clk game.writer.tracker.next_frame\[295\] net1281 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[295\] sky130_fd_sc_hd__dfrtp_1
X_12035_ _05235_ _05237_ _05240_ _05242_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__or4_1
X_17892_ net615 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_256_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19631_ clknet_leaf_28_clk game.writer.tracker.next_frame\[226\] net1309 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[226\] sky130_fd_sc_hd__dfrtp_1
X_16843_ net132 net53 net142 _02617_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[236\]
+ sky130_fd_sc_hd__a31o_1
XANTENNA__16615__A2 _02524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14211__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_189_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19562_ clknet_leaf_37_clk game.writer.tracker.next_frame\[157\] net1349 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[157\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16774_ _02435_ net64 _02593_ net1938 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[191\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12012__A _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15026__C net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13986_ net942 game.CPU.applesa.ab.check_walls.above.walls\[23\] vssd1 vssd1 vccd1
+ vccd1 _07860_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_358_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18513_ net579 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__inv_2
XANTENNA__09502__B1 game.CPU.applesa.ab.check_walls.above.walls\[51\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_358_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15725_ game.CPU.applesa.ab.absxs.body_x\[53\] net473 vssd1 vssd1 vccd1 vccd1 _01737_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output35_A net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12937_ _06720_ _06721_ net688 vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__mux2_1
X_19493_ clknet_leaf_24_clk game.writer.tracker.next_frame\[88\] net1338 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[88\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10112__A1 game.CPU.applesa.enable_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09799__Y _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_272_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17040__A2 _02678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18444_ net592 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_272_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10663__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15656_ game.CPU.applesa.ab.check_walls.above.walls\[52\] net342 vssd1 vssd1 vccd1
+ vccd1 _01668_ sky130_fd_sc_hd__nand2_1
X_12868_ game.writer.tracker.frame\[290\] game.writer.tracker.frame\[291\] net988
+ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_199_Right_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14607_ game.CPU.clock1.counter\[7\] _08460_ net267 vssd1 vssd1 vccd1 vccd1 _08462_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18375_ net597 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15042__B net1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11819_ game.CPU.applesa.ab.check_walls.above.walls\[29\] net308 _05706_ vssd1 vssd1
+ vccd1 vccd1 _05707_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09805__A1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10467__A game.CPU.applesa.ab.absxs.body_x\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15587_ _03396_ net356 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__nand2_1
X_12799_ _06669_ _06670_ _06672_ _06671_ net493 net691 vssd1 vssd1 vccd1 vccd1 _06673_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09805__B2 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17326_ net130 _02592_ net732 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14538_ _08406_ _08408_ vssd1 vssd1 vccd1 vccd1 _08411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16000__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17257_ net111 _02467_ _02745_ net1935 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[522\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_330_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16551__A1 _02237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14469_ game.CPU.applesa.ab.absxs.body_x\[62\] net1058 vssd1 vssd1 vccd1 vccd1 _08343_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__12682__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13365__A1 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16208_ _02020_ _02021_ _02024_ _02025_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__or4_1
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12799__S0 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_231_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17188_ _02494_ net71 net727 vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__o21a_1
XFILLER_0_302_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16139_ _02084_ _02088_ _02091_ _02070_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__o31a_1
XANTENNA__15993__A game.CPU.applesa.ab.check_walls.above.walls\[98\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16854__A2 _02623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08961_ game.CPU.apple_location\[0\] vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__inv_2
XANTENNA__13668__A2 _07541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_282_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17803__A1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19829_ clknet_leaf_38_clk game.writer.tracker.next_frame\[424\] net1329 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[424\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_320_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_235_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18996__CLK net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12628__B1 game.CPU.applesa.twoapples.absxs.next_head\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_242_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13825__C1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14093__A2 game.CPU.applesa.ab.check_walls.above.walls\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09513_ net1093 _03272_ _03273_ net1111 vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__o22a_1
XFILLER_0_149_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16329__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10103__B2 _04256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11300__B1 _05189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13840__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19350__D game.CPU.applesa.twoapples.absxs.next_head\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_A _08416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17031__A2 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11761__A game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ net1126 game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1 vssd1 vccd1
+ vccd1 _03687_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_84_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11851__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11480__B net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_325_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ net1086 game.CPU.applesa.ab.check_walls.above.walls\[11\] vssd1 vssd1 vccd1
+ vccd1 _03618_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10377__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16790__A1 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout523_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15593__A2 game.CPU.walls.rand_wall.abduyd.next_wall\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1265_A game.CPU.applesa.ab.absxs.body_x\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15887__B net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_331_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19621__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09885__B _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__X _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1053_X net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_144_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout892_A net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17098__A2 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16214__D _02225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1220_X net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13108__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10150_ game.CPU.randy.f1.state\[2\] game.CPU.randy.f1.state\[1\] game.CPU.randy.f1.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__or3b_1
XANTENNA__19771__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18987__Q game.CPU.applesa.ab.check_walls.above.walls\[32\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17607__B net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13627__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11936__A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10081_ _04219_ _04220_ net1153 vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_167_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_261_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_342_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_273_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09406__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19001__CLK net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout945_X net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12528__A2_N net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17270__A2 _02327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ game.writer.tracker.frame\[523\] net708 net671 game.writer.tracker.frame\[524\]
+ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__o22a_1
XANTENNA__10893__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13771_ game.writer.tracker.frame\[159\] net711 net674 game.writer.tracker.frame\[160\]
+ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__o22a_1
X_10983_ _04866_ _04867_ _04871_ _04872_ _04870_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a221o_1
XANTENNA__13362__S net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13831__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16239__A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15510_ _01532_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__inv_2
XANTENNA__15143__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ _06571_ _06593_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16490_ game.writer.tracker.frame\[64\] _02433_ _02436_ _02273_ vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[64\] sky130_fd_sc_hd__a22o_1
XANTENNA__11842__A1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_247_Left_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12486__B net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09141__A game.CPU.applesa.ab.check_walls.above.walls\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15441_ _08917_ _08931_ _01467_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_194_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18719__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12653_ game.CPU.applesa.ab.absxs.body_x\[7\] net531 net360 game.CPU.applesa.ab.absxs.body_y\[4\]
+ _06245_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__o221a_1
XANTENNA__16781__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14982__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_178_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11799__A2_N net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11604_ net779 _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__xnor2_1
X_18160_ net630 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__inv_2
X_15372_ _08904_ _08913_ vssd1 vssd1 vccd1 vccd1 _08914_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15797__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_191_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ _03291_ game.CPU.applesa.twoapples.absxs.next_head\[1\] net372 game.CPU.applesa.ab.absxs.body_x\[10\]
+ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__a22o_1
X_17111_ net161 net56 net81 _02705_ net1469 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[416\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14323_ game.CPU.applesa.ab.absxs.body_x\[75\] net1046 vssd1 vssd1 vccd1 vccd1 _08197_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_312_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18091_ net589 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__inv_2
X_11535_ net790 net249 vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__and2_1
XANTENNA__11070__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16533__A1 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17042_ _02535_ _02670_ net726 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__o21a_1
XANTENNA__14544__B1 _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_311_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14254_ _08119_ _08120_ _08126_ _08127_ vssd1 vssd1 vccd1 vccd1 _08128_ sky130_fd_sc_hd__a22o_1
X_11466_ game.CPU.applesa.ab.check_walls.above.walls\[16\] net777 vssd1 vssd1 vccd1
+ vccd1 _05355_ sky130_fd_sc_hd__xnor2_1
X_13205_ game.writer.tracker.frame\[428\] game.writer.tracker.frame\[429\] net1020
+ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__mux2_1
X_10417_ _04359_ _04562_ _04561_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_256_Left_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11397_ game.CPU.applesa.ab.check_walls.above.walls\[88\] net778 vssd1 vssd1 vccd1
+ vccd1 _05286_ sky130_fd_sc_hd__xnor2_1
X_14185_ _03354_ net987 net860 game.CPU.applesa.ab.absxs.body_y\[19\] _08058_ vssd1
+ vssd1 vccd1 vccd1 _08059_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_267_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16836__A2 _02375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ game.writer.tracker.frame\[166\] game.writer.tracker.frame\[167\] net990
+ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__mux2_1
XANTENNA__09971__B1 _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10348_ game.CPU.walls.rand_wall.counter2\[2\] game.CPU.walls.rand_wall.counter2\[1\]
+ game.CPU.walls.rand_wall.counter2\[0\] vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_209_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ net1197 _00219_ _00664_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_280_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13067_ game.writer.tracker.frame\[214\] game.writer.tracker.frame\[215\] net1027
+ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17944_ net655 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__inv_2
X_10279_ net1166 _04257_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_268_Right_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_252_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09316__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11565__B net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ game.CPU.applesa.ab.check_walls.above.walls\[44\] net554 vssd1 vssd1 vccd1
+ vccd1 _05905_ sky130_fd_sc_hd__or2_1
X_17875_ net636 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__inv_2
XFILLER_0_233_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19614_ clknet_leaf_27_clk game.writer.tracker.next_frame\[209\] net1310 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[209\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17261__A2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16826_ net131 _02609_ _02607_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[227\]
+ sky130_fd_sc_hd__a21o_1
XANTENNA__12038__A1_N game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16757_ _02405_ net100 net736 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__o21a_1
X_19545_ clknet_leaf_49_clk game.writer.tracker.next_frame\[140\] net1297 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[140\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_265_Left_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13969_ net1045 game.CPU.applesa.ab.check_walls.above.walls\[83\] vssd1 vssd1 vccd1
+ vccd1 _07843_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_232_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12677__A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19170__D _00288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17013__A2 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15708_ _03461_ net336 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_278_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19476_ clknet_leaf_19_clk game.writer.tracker.next_frame\[71\] net1335 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[71\] sky130_fd_sc_hd__dfrtp_1
X_16688_ net204 net68 net62 _02563_ net1770 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[135\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_291_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09051__A game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_173_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15639_ game.CPU.applesa.ab.absxs.body_y\[80\] net449 vssd1 vssd1 vccd1 vccd1 _01651_
+ sky130_fd_sc_hd__xnor2_1
X_18427_ net588 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16772__A1 _02429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19644__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_347_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_302_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09160_ game.CPU.applesa.ab.check_walls.above.walls\[53\] vssd1 vssd1 vccd1 vccd1
+ _03409_ sky130_fd_sc_hd__inv_2
X_18358_ net596 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17309_ net1989 net723 _02759_ _02397_ net176 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[560\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_83_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15500__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09091_ game.CPU.applesa.ab.absxs.body_y\[56\] vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__inv_2
XFILLER_0_161_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16524__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18289_ net618 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_342_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19794__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_274_Left_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_287_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload43_A clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14116__B net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13433__S1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_330_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout104_A net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16827__A2 _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13955__B net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ game.CPU.apple_location\[6\] game.CPU.applesa.ab.apple_location\[6\] _04207_
+ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_244_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08944_ net1101 vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__inv_2
XANTENNA__14132__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1013_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13510__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09226__A game.CPU.applesa.ab.check_walls.above.walls\[176\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_235_Right_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20001__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__B net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout473_A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18539__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13971__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17252__A2 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19174__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_283_Left_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16460__B1 _02416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout640_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout738_A _04738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11491__A game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_338_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09427_ net1098 game.CPU.applesa.ab.check_walls.above.walls\[113\] vssd1 vssd1 vccd1
+ vccd1 _03670_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16763__A1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1170_X net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09358_ net1088 game.CPU.applesa.ab.check_walls.above.walls\[195\] vssd1 vssd1 vccd1
+ vccd1 _03601_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11815__A1_N net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16515__A1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09289_ net1137 net809 vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__or2_1
XFILLER_0_306_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_292_Left_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13329__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11320_ game.CPU.applesa.ab.apple_possible\[4\] _04462_ vssd1 vssd1 vccd1 vccd1 _05209_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10260__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ game.CPU.applesa.ab.absxs.body_x\[114\] net409 net545 game.CPU.applesa.ab.absxs.body_x\[115\]
+ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_344_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10202_ net1089 _04394_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16818__A2 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11182_ game.CPU.applesa.ab.absxs.body_y\[85\] net543 vssd1 vssd1 vccd1 vccd1 _05072_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_293_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11666__A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ game.CPU.randy.f1.c1.max_i\[0\] game.CPU.randy.f1.c1.count\[0\] vssd1 vssd1
+ vccd1 vccd1 _04328_ sky130_fd_sc_hd__xor2_1
XANTENNA__15138__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14042__A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15990_ _01994_ _01995_ _01996_ _02001_ _01989_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__o41a_1
XANTENNA__17491__A2 _02778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19517__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_234_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13501__A1 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _04268_ _04271_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__xnor2_1
X_14941_ _08714_ _08717_ vssd1 vssd1 vccd1 vccd1 _08718_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09136__A game.CPU.applesa.ab.check_walls.above.walls\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_202_Right_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18449__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17243__A2 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17660_ _03052_ net194 _03051_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__and3b_1
XFILLER_0_199_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14872_ game.CPU.walls.abc.number\[4\] game.CPU.walls.abc.number\[0\] game.CPU.walls.abc.counter
+ vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__mux2_1
X_16611_ net177 _02480_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_106_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13823_ net285 _07688_ _07695_ _07696_ net242 vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__a221o_1
XFILLER_0_202_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17591_ _03009_ _03010_ net582 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__a21oi_1
XANTENNA__19667__CLK clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_355_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13804__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16542_ net202 net146 _02310_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__and3_1
X_19330_ clknet_leaf_72_clk net1413 _00935_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twomode.number\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_13754_ game.writer.tracker.frame\[165\] game.writer.tracker.frame\[167\] game.writer.tracker.frame\[168\]
+ game.writer.tracker.frame\[166\] net969 net990 vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11815__B2 _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10966_ net1265 net406 vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ _06554_ _06564_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__nand2_1
X_19261_ clknet_leaf_8_clk _00049_ _00891_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count1\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_16473_ net1882 _02420_ _02424_ net112 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[59\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16754__A1 _02398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12784__X _06658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13685_ game.writer.tracker.frame\[485\] game.writer.tracker.frame\[487\] game.writer.tracker.frame\[488\]
+ game.writer.tracker.frame\[486\] net974 net999 vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__mux4_1
XANTENNA__11291__A2 _04949_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10897_ game.CPU.applesa.ab.check_walls.collision_up _04797_ vssd1 vssd1 vccd1 vccd1
+ _04799_ sky130_fd_sc_hd__and2_1
XANTENNA__13820__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18212_ net664 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__inv_2
X_15424_ net833 _01444_ _08935_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15601__A game.CPU.applesa.ab.check_walls.above.walls\[112\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_344_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19192_ clknet_leaf_46_clk net345 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.x_final\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_12636_ _06393_ _06395_ _06396_ _06397_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18691__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_316_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18143_ net630 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__inv_2
XFILLER_0_344_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15355_ _08887_ _08896_ _08894_ vssd1 vssd1 vccd1 vccd1 _08897_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_5_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12567_ game.CPU.applesa.ab.absxs.body_x\[117\] net378 game.CPU.applesa.twoapples.absxs.next_head\[4\]
+ _03355_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ game.CPU.applesa.ab.absxs.body_x\[28\] net1070 vssd1 vssd1 vccd1 vccd1 _08180_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_215_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18074_ net657 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__inv_2
X_11518_ _03380_ net256 vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__xnor2_1
X_15286_ _01264_ _08817_ _08818_ _08827_ _01265_ vssd1 vssd1 vccd1 vccd1 _08838_ sky130_fd_sc_hd__a41o_1
XPHY_EDGE_ROW_337_Right_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_269_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12498_ game.CPU.applesa.ab.absxs.body_x\[64\] net382 vssd1 vssd1 vccd1 vccd1 _06375_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19047__CLK net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold208 game.writer.tracker.frame\[365\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
X_17025_ _02521_ _02663_ _02677_ net1680 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[356\]
+ sky130_fd_sc_hd__a22o_1
Xhold219 game.writer.tracker.frame\[527\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14237_ _08107_ _08108_ _08109_ _08110_ vssd1 vssd1 vccd1 vccd1 _08111_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11449_ game.CPU.applesa.ab.check_walls.above.walls\[75\] net763 vssd1 vssd1 vccd1
+ vccd1 _05338_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16809__A2 _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14168_ game.CPU.applesa.ab.absxs.body_y\[104\] net989 vssd1 vssd1 vccd1 vccd1 _08042_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_237_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10554__B2 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13267__S net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13119_ game.writer.tracker.frame\[170\] game.writer.tracker.frame\[171\] net990
+ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15048__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10480__A _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14099_ _07963_ _07965_ _07967_ _07972_ vssd1 vssd1 vccd1 vccd1 _07973_ sky130_fd_sc_hd__or4_4
X_18976_ net1196 _00201_ _00647_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_252_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09046__A game.CPU.applesa.ab.absxs.body_y\[100\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17927_ net613 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__inv_2
XANTENNA__14887__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1270 game.CPU.applesa.ab.absxs.body_y\[63\] vssd1 vssd1 vccd1 vccd1 net1270
+ sky130_fd_sc_hd__buf_2
XANTENNA__17234__A2 _02422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1281 net1360 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__clkbuf_4
Xfanout1292 net1293 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__buf_2
X_17858_ _03180_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__inv_2
XFILLER_0_205_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_233_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16809_ net150 _02497_ net104 _02603_ net1822 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[216\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_220_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17789_ _01263_ _08818_ _08827_ _01264_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a31o_1
XANTENNA__15796__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19528_ clknet_leaf_23_clk game.writer.tracker.next_frame\[123\] net1347 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[123\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10609__A2 _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12200__A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_354_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19459_ clknet_leaf_39_clk game.writer.tracker.next_frame\[54\] net1352 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[54\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_313_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13559__A1 game.writer.tracker.frame\[98\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09212_ game.CPU.applesa.ab.check_walls.above.walls\[157\] vssd1 vssd1 vccd1 vccd1
+ _03461_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14220__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13654__S1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09143_ game.CPU.applesa.ab.check_walls.above.walls\[26\] vssd1 vssd1 vccd1 vccd1
+ _03392_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13669__C _07504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_A game.CPU.applesa.ab.absxs.next_head\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09074_ game.CPU.applesa.ab.absxs.body_y\[113\] vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__inv_2
XFILLER_0_288_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17170__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_250_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_304_Right_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1130_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout107_X net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1228_A game.CPU.walls.rand_wall.start_enable vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19565__RESET_B net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_275_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout590_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16061__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_338_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09976_ net1148 net848 _04203_ vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__a21o_1
XANTENNA__15484__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14287__A2 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15484__B2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18564__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13590__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17225__A2 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_354_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11933__B net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16984__A1 _02465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19161__Q game.CPU.walls.rand_wall.input2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13342__S0 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10820_ game.CPU.applesa.ab.absxs.body_y\[9\] _04689_ _04707_ game.CPU.applesa.ab.absxs.body_y\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__a22o_1
XANTENNA__17901__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_357_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10751_ game.CPU.applesa.ab.absxs.body_y\[112\] _04663_ _04664_ game.CPU.applesa.ab.absxs.body_y\[108\]
+ vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__a22o_1
XANTENNA__12470__A1 game.CPU.applesa.ab.absxs.body_x\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_149_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16736__A1 net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12470__B2 game.CPU.applesa.ab.absxs.body_y\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_223_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout908_X net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_326_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13470_ net704 _07084_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_175_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10682_ game.CPU.applesa.ab.absxs.body_x\[10\] _04689_ _04707_ game.CPU.applesa.ab.absxs.body_x\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_350_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16236__B net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ game.CPU.applesa.ab.absxs.body_x\[33\] net375 net529 game.CPU.applesa.ab.absxs.body_x\[35\]
+ _06296_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__o221a_1
XFILLER_0_326_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15140__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15140_ net1210 net1236 game.CPU.applesa.ab.check_walls.above.walls\[168\] vssd1
+ vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__and3_1
XANTENNA__13970__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12352_ game.CPU.applesa.ab.absxs.body_y\[79\] net367 vssd1 vssd1 vccd1 vccd1 _06229_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__17161__A1 _02450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13970__B2 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16523__Y _02462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10784__B2 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11303_ game.CPU.applesa.ab.apple_possible\[5\] _04775_ vssd1 vssd1 vccd1 vccd1 _05192_
+ sky130_fd_sc_hd__or2_2
X_15071_ net1217 net1246 game.CPU.applesa.ab.check_walls.above.walls\[99\] vssd1 vssd1
+ vccd1 vccd1 _00096_ sky130_fd_sc_hd__and3_1
X_12283_ _06035_ _06168_ _06037_ _06036_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_294_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_189_Left_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14022_ net881 game.CPU.applesa.ab.check_walls.above.walls\[161\] vssd1 vssd1 vccd1
+ vccd1 _07896_ sky130_fd_sc_hd__nor2_1
XANTENNA__09926__B1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ game.CPU.applesa.ab.absxs.body_y\[14\] net539 vssd1 vssd1 vccd1 vccd1 _05124_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__17067__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10536__A1 game.CPU.applesa.ab.absxs.body_x\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_264_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18907__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18830_ clknet_leaf_3_clk _01221_ _00558_ vssd1 vssd1 vccd1 vccd1 game.CPU.bodymain1.Direction\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_11165_ game.CPU.applesa.ab.absxs.body_y\[50\] net538 net416 game.CPU.applesa.ab.absxs.body_x\[48\]
+ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_248_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15475__A1 _01454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ game.CPU.applesa.enable_in game.CPU.applesa.twoapples.x_final\[2\] _03212_
+ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__a21o_1
X_11096_ game.CPU.applesa.ab.absxs.body_x\[56\] net415 vssd1 vssd1 vccd1 vccd1 _04986_
+ sky130_fd_sc_hd__xnor2_1
X_15973_ _03269_ net356 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__nand2_1
X_18761_ clknet_leaf_12_clk _01178_ _00498_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[55\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_207_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_303_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10047_ net1274 net1271 vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__nor2_1
X_17712_ net1271 _04435_ _03083_ _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__o211a_2
X_14924_ _08697_ _08700_ vssd1 vssd1 vccd1 vccd1 _08701_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13581__S0 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap66_A _02514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18692_ clknet_leaf_58_clk _01109_ _00429_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[34\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold80 game.writer.tracker.frame\[438\] vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_264_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold91 net43 vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_349_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14004__A1_N net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17643_ _08803_ net194 _03041_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__and3_1
X_14855_ game.CPU.randy.f1.c1.count\[10\] _08645_ net2023 vssd1 vssd1 vccd1 vccd1
+ _08648_ sky130_fd_sc_hd__a21oi_1
XANTENNA__16975__A1 net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13806_ net495 _07677_ _07678_ _07679_ net215 vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__a311o_1
XPHY_EDGE_ROW_198_Left_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17574_ net1259 _02843_ _02854_ _02997_ _02830_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__a2111o_1
X_14786_ _08604_ vssd1 vssd1 vccd1 vccd1 _08605_ sky130_fd_sc_hd__inv_2
XANTENNA__15034__C game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_201_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11998_ _05882_ _05883_ _05884_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_67_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16525_ net167 _02286_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_275_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19313_ net1164 _00037_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.out_random_2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13737_ game.writer.tracker.frame\[213\] game.writer.tracker.frame\[215\] game.writer.tracker.frame\[216\]
+ game.writer.tracker.frame\[214\] net978 net1027 vssd1 vssd1 vccd1 vccd1 _07611_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_280_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10949_ game.CPU.applesa.ab.absxs.body_x\[30\] net411 net396 game.CPU.applesa.ab.absxs.body_y\[31\]
+ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__a22o_1
XANTENNA__11264__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12955__A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_217_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_70_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_8
X_16456_ net171 _02328_ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__or2_4
X_19244_ clknet_leaf_17_clk _00058_ _00882_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_280_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13668_ _07540_ _07541_ net179 vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16146__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15407_ _01432_ _01434_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15050__B net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19175_ clknet_leaf_4_clk _01294_ _00837_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12619_ net1267 net384 _06228_ _06486_ _06495_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__a2111o_1
X_16387_ net189 net205 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__nor2_1
X_13599_ game.writer.tracker.frame\[301\] game.writer.tracker.frame\[303\] game.writer.tracker.frame\[304\]
+ game.writer.tracker.frame\[302\] net964 net989 vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18126_ net577 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__inv_2
XFILLER_0_289_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15338_ game.writer.updater.commands.cmd_num\[1\] game.writer.updater.commands.cmd_num\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08880_ sky130_fd_sc_hd__xor2_1
XFILLER_0_206_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17152__A1 _02429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15985__B net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13961__B2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16433__Y _02396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18057_ net629 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__inv_2
X_15269_ _08819_ _08820_ _08824_ vssd1 vssd1 vccd1 vccd1 _08825_ sky130_fd_sc_hd__or3_1
XFILLER_0_340_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17008_ _02494_ _02638_ net728 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_286_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10527__A1 game.CPU.applesa.ab.absxs.body_x\[55\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18587__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__B2 game.CPU.applesa.ab.absxs.body_x\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09393__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout507 net516 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_228_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ net1132 _03318_ _03319_ net1149 _04066_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19832__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16258__A3 _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09393__B2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout518 _06214_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_2
Xfanout529 net532 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14269__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09761_ net1112 _03390_ _03394_ net1150 _04003_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__a221o_1
X_18959_ net1201 _00232_ _00630_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17207__A2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13572__S0 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_280_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09692_ net1100 game.CPU.applesa.ab.absxs.body_x\[5\] vssd1 vssd1 vccd1 vccd1 _03935_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16415__B1 _02383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09696__A2 game.CPU.applesa.ab.absxs.body_y\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19982__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16140__A1_N net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13229__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16966__A1 _02428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout171_A net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13324__S0 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_A game.CPU.walls.rand_wall.abduyd.next_wall\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_317_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16430__A3 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_239_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11255__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1080_A game.CPU.bad_collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_61_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout436_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1178_A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout224_X net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1345_A net1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09126_ net965 vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__inv_2
XFILLER_0_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19362__CLK clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15895__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17143__A1 net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16343__Y _02331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__A2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10766__B2 game.CPU.applesa.ab.absxs.body_y\[78\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_161_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09057_ game.CPU.applesa.ab.absxs.body_y\[54\] vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__inv_2
XANTENNA__09893__B _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_328_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_248_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1133_X net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_276_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold550 game.writer.tracker.frame\[522\] vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 game.writer.tracker.frame\[534\] vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout972_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold572 game.writer.tracker.frame\[469\] vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11715__B1 game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold583 game.writer.tracker.frame\[552\] vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_291_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09384__B2 net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17446__A2 _02779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 game.writer.tracker.frame\[31\] vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout84_A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _04187_ _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ _06655_ _06656_ net682 vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11663__B net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09414__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _05793_ _05794_ _05799_ _05808_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__o31a_1
XANTENNA__16957__A1 _02412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_339_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ net1985 _08480_ _08482_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[19\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_358_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11852_ net819 net302 _05735_ _05736_ _05739_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_352_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10279__B _04257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14432__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_358_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10803_ game.CPU.applesa.ab.absxs.body_y\[26\] _04695_ _04698_ game.CPU.applesa.ab.absxs.body_y\[22\]
+ vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14571_ net929 _08432_ vssd1 vssd1 vccd1 vccd1 _08434_ sky130_fd_sc_hd__nand2_1
XANTENNA__11246__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16709__A1 _02238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_220_Left_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11783_ _05664_ _05669_ _05670_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_52_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13370__S net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16310_ _02283_ _02306_ _02305_ _08028_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a2bb2o_1
X_13522_ net247 _07394_ _07395_ _07341_ net191 vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__a221o_1
XANTENNA__15151__A net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17290_ net116 net156 net66 _02754_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[546\]
+ sky130_fd_sc_hd__a31o_1
X_10734_ game.CPU.applesa.ab.absxs.body_y\[21\] _04645_ _04652_ game.CPU.applesa.ab.absxs.body_y\[17\]
+ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__a22o_1
XANTENNA__19705__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16185__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16241_ _06607_ _02226_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__and2b_1
XFILLER_0_353_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13453_ _07023_ _07028_ net705 vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_341_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10665_ net1080 _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nor2_2
XFILLER_0_326_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16534__X _02470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13943__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12404_ game.CPU.applesa.ab.absxs.body_x\[52\] net382 vssd1 vssd1 vccd1 vccd1 _06281_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_341_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16172_ game.CPU.applesa.ab.absxs.body_x\[33\] net472 net451 game.CPU.applesa.ab.absxs.body_y\[32\]
+ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a22o_1
XANTENNA__17134__A1 _02394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13384_ _06863_ _06881_ net680 vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__mux2_1
XANTENNA__13943__B2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17349__Y _02779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ game.CPU.applesa.ab.absxs.body_x\[98\] net263 _04669_ net929 vssd1 vssd1
+ vccd1 vccd1 _01141_ sky130_fd_sc_hd__a22o_1
XANTENNA__19416__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15123_ net1207 net1230 net789 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_212_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12335_ net517 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.absxs.next_head\[6\]
+ sky130_fd_sc_hd__clkinv_4
XANTENNA__19855__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_322_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_188_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13156__C1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19931_ clknet_leaf_48_clk game.writer.tracker.next_frame\[526\] net1302 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[526\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16893__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15054_ net1218 net1247 game.CPU.applesa.ab.check_walls.above.walls\[82\] vssd1 vssd1
+ vccd1 vccd1 _00277_ sky130_fd_sc_hd__and3_1
XFILLER_0_294_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12266_ game.CPU.applesa.ab.check_walls.above.walls\[109\] net548 vssd1 vssd1 vccd1
+ vccd1 _06152_ sky130_fd_sc_hd__nand2_1
XANTENNA__10742__B _04658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14005_ net867 game.CPU.applesa.ab.check_walls.above.walls\[140\] net791 net852 _07876_
+ vssd1 vssd1 vccd1 vccd1 _07879_ sky130_fd_sc_hd__a221o_1
X_11217_ _03244_ net410 vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__nand2_1
X_19862_ clknet_leaf_20_clk game.writer.tracker.next_frame\[457\] net1315 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[457\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09308__B game.CPU.applesa.ab.absxs.body_x\[53\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_281_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12197_ net818 net423 vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_247_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18813_ clknet_leaf_72_clk game.CPU.clock1.next_counter\[16\] _00550_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_247_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11148_ game.CPU.applesa.ab.absxs.body_x\[99\] net408 vssd1 vssd1 vccd1 vccd1 _05038_
+ sky130_fd_sc_hd__nand2_1
X_19793_ clknet_leaf_35_clk game.writer.tracker.next_frame\[388\] net1355 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[388\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15999__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13545__S net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13554__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18744_ clknet_leaf_11_clk _01161_ _00481_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16660__A3 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15956_ game.CPU.applesa.ab.check_walls.above.walls\[28\] net453 vssd1 vssd1 vccd1
+ vccd1 _01968_ sky130_fd_sc_hd__xnor2_1
X_11079_ game.CPU.applesa.ab.absxs.body_x\[43\] net544 net538 game.CPU.applesa.ab.absxs.body_y\[42\]
+ _04965_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__o221a_1
XANTENNA__12131__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09678__A2 game.CPU.applesa.ab.absxs.body_y\[103\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_223_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14907_ _08669_ _08677_ _08680_ _08683_ vssd1 vssd1 vccd1 vccd1 _08684_ sky130_fd_sc_hd__and4_1
XANTENNA__16948__A1 _02394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19235__CLK clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15887_ game.CPU.applesa.ab.check_walls.above.walls\[140\] net450 vssd1 vssd1 vccd1
+ vccd1 _01899_ sky130_fd_sc_hd__xnor2_1
X_18675_ clknet_leaf_8_clk _01092_ _00412_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_349_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_199_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17070__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17626_ _03032_ net429 _03031_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__and3b_1
XFILLER_0_156_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14838_ _04327_ _08633_ _08637_ _04332_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[4\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_187_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14423__A2 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_203_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12434__A1 net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14769_ _08587_ _08588_ _08589_ vssd1 vssd1 vccd1 vccd1 _08590_ sky130_fd_sc_hd__or3_1
X_17557_ net739 _02851_ _02951_ _02845_ _02982_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__a221o_1
XANTENNA__13631__B1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12685__A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_336_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_323_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16508_ net219 _02362_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__nor2_8
XANTENNA__19385__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17488_ net1121 _04628_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_9_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19227_ clknet_leaf_57_clk _00020_ _00865_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.normal1.number\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_15_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16439_ net1278 _07916_ _08027_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__or3b_4
XANTENNA__14187__B2 game.CPU.applesa.ab.absxs.body_y\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_344_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18372__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_288_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13395__C1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13934__A1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17125__A1 _02379_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19158_ clknet_leaf_3_clk _01279_ _00829_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.counter2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13934__B2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16604__B _02480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18109_ net632 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__inv_2
XANTENNA__10933__A game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19089_ net1178 _00126_ _00760_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[134\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_258_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_257_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_300_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_285_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14124__B game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_273_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_319_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout304 _05608_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_238_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16620__A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout315 _05213_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_4
X_20002_ clknet_leaf_44_clk game.writer.updater.update.next\[0\] net1300 vssd1 vssd1
+ vccd1 vccd1 game.writer.updater.commands.mode\[0\] sky130_fd_sc_hd__dfrtp_4
Xfanout326 game.CPU.applesa.ab.absxs.next_head\[0\] vssd1 vssd1 vccd1 vccd1 net326
+ sky130_fd_sc_hd__clkbuf_8
Xfanout337 net340 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_8
X_09813_ net911 game.CPU.applesa.ab.absxs.body_x\[24\] game.CPU.applesa.ab.absxs.body_y\[27\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__a22o_1
Xfanout348 net349 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_4
Xfanout359 net363 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_323_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout386_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ net1131 game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1 vccd1
+ vccd1 _03987_ sky130_fd_sc_hd__xor2_1
XFILLER_0_185_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_161_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12579__B net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ net1085 net1265 vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout174_X net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16939__A1 net148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1295_A net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19728__CLK clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18602__CLK clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14414__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19998__RESET_B net1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13622__A0 game.writer.tracker.frame\[273\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout720_A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_34_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_X net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A game.CPU.applesa.ab.check_walls.above.walls\[55\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10436__B1 _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16167__A2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18752__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19878__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18282__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1348_X net1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10450_ _04582_ _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__and2_1
XFILLER_0_323_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17116__A1 _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10739__A1 game.CPU.applesa.ab.absxs.body_y\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10739__B2 game.CPU.applesa.ab.absxs.body_y\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09109_ net1460 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__inv_2
X_10381_ net919 game.CPU.apple_location2\[2\] game.CPU.apple_location2\[6\] net902
+ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_115_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12120_ game.CPU.applesa.ab.check_walls.above.walls\[172\] net552 vssd1 vssd1 vccd1
+ vccd1 _06007_ sky130_fd_sc_hd__or2_1
XANTENNA__09409__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout975_X net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14034__B game.CPU.applesa.ab.check_walls.above.walls\[112\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09357__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09357__B2 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ game.CPU.applesa.ab.check_walls.above.walls\[61\] net389 vssd1 vssd1 vccd1
+ vccd1 _05938_ sky130_fd_sc_hd__xnor2_1
Xhold380 game.writer.tracker.frame\[516\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold391 game.writer.tracker.frame\[468\] vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_263_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11164__A1 game.CPU.applesa.ab.absxs.body_y\[50\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_261_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11002_ game.CPU.applesa.ab.absxs.body_x\[47\] net545 net539 game.CPU.applesa.ab.absxs.body_y\[46\]
+ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a22o_1
XANTENNA__19614__Q game.writer.tracker.frame\[209\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_183_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout860 _03376_ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_4
XANTENNA__11674__A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13536__S0 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout871 net872 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_4
XANTENNA__15146__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15810_ _03414_ net338 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__xnor2_1
X_16790_ net147 _02467_ net102 _02598_ net1487 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[202\]
+ sky130_fd_sc_hd__a32o_1
Xfanout882 net885 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_125_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout893 net895 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_300_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12489__B net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09144__A game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15741_ _03474_ game.CPU.walls.rand_wall.abduyd.next_wall\[7\] vssd1 vssd1 vccd1
+ vccd1 _01753_ sky130_fd_sc_hd__nor2_1
XANTENNA__11393__B net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ net205 _06751_ _06826_ net281 vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__a211o_1
XANTENNA__14985__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11904_ game.CPU.applesa.ab.check_walls.above.walls\[92\] net393 net302 game.CPU.applesa.ab.check_walls.above.walls\[94\]
+ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__o22a_1
XFILLER_0_169_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15672_ game.CPU.applesa.ab.check_walls.above.walls\[10\] net348 vssd1 vssd1 vccd1
+ vccd1 _01684_ sky130_fd_sc_hd__nand2_1
X_18460_ net654 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__inv_2
X_12884_ game.writer.tracker.frame\[12\] game.writer.tracker.frame\[13\] net1004 vssd1
+ vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_358_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09431__X _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_319_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14623_ game.CPU.clock1.counter\[13\] _08470_ net267 vssd1 vssd1 vccd1 vccd1 _08472_
+ sky130_fd_sc_hd__o21ai_1
X_17411_ net1275 _02840_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__or2_2
XFILLER_0_185_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11835_ net790 net390 net299 game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1
+ vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__o2bb2a_1
X_18391_ net599 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_2
XANTENNA__13613__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_25_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_272_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_346_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17342_ game.CPU.kyle.L1.nextState\[5\] game.CPU.kyle.L1.nextState\[4\] vssd1 vssd1
+ vccd1 vccd1 _02772_ sky130_fd_sc_hd__nor2_2
XFILLER_0_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14554_ game.CPU.walls.rand_wall.logic_enable _08421_ _08422_ vssd1 vssd1 vccd1 vccd1
+ _08423_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11766_ game.CPU.applesa.ab.check_walls.above.walls\[182\] net301 _05648_ _05649_
+ _05653_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14209__B net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13505_ net247 _07375_ _07377_ _07378_ _07326_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__o32a_1
X_17273_ _02278_ _02491_ _02749_ net1946 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[534\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_194_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10717_ game.CPU.applesa.ab.absxs.body_y\[53\] _04609_ _04637_ game.CPU.applesa.ab.absxs.body_y\[49\]
+ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14485_ _08319_ _08320_ _08323_ _08072_ vssd1 vssd1 vccd1 vccd1 _08359_ sky130_fd_sc_hd__o31a_2
XFILLER_0_138_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16264__X _02270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11697_ game.CPU.applesa.ab.check_walls.above.walls\[160\] net774 vssd1 vssd1 vccd1
+ vccd1 _05586_ sky130_fd_sc_hd__xor2_1
XFILLER_0_43_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13377__C1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16224_ _08028_ net141 _02232_ net1932 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[2\]
+ sky130_fd_sc_hd__a22o_1
X_19012_ net1196 _00240_ _00683_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[57\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_341_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13436_ _07308_ _07309_ net491 vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17107__A1 net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10648_ game.CPU.bad_collision _03245_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__nor2_1
XANTENNA__16424__B _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_341_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16155_ _01716_ _02166_ _01720_ _02165_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__or4b_2
XANTENNA__11849__A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13367_ net278 _07234_ _07239_ _07240_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__o22a_1
X_10579_ net936 game.CPU.applesa.ab.absxs.body_x\[100\] _04657_ _04662_ vssd1 vssd1
+ vccd1 vccd1 _01151_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15106_ net1205 net1232 game.CPU.applesa.ab.check_walls.above.walls\[134\] vssd1
+ vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__and3_1
XANTENNA__16866__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12318_ _06199_ _06200_ _06201_ _06203_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__and4_1
XANTENNA__11568__B net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16086_ game.CPU.applesa.ab.check_walls.above.walls\[150\] net439 net430 net789 vssd1
+ vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__a2bb2o_1
X_13298_ net513 _07169_ _07171_ net215 vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19914_ clknet_leaf_23_clk game.writer.tracker.next_frame\[509\] net1344 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[509\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_286_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_283_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15037_ net1219 net1245 game.CPU.applesa.ab.check_walls.above.walls\[65\] vssd1 vssd1
+ vccd1 vccd1 _00258_ sky130_fd_sc_hd__and3_1
X_12249_ _05988_ _05989_ _06133_ _06134_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__or4_2
XFILLER_0_294_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_282_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_225_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_299_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_286_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19845_ clknet_leaf_36_clk game.writer.tracker.next_frame\[440\] net1357 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[440\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_273_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17267__A2_N _02403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15056__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19776_ clknet_leaf_26_clk game.writer.tracker.next_frame\[371\] net1312 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[371\] sky130_fd_sc_hd__dfrtp_1
X_16988_ _02470_ net88 _02667_ net1500 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[331\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12104__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18625__CLK clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12399__B net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18727_ clknet_leaf_13_clk _01144_ _00464_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[109\]
+ sky130_fd_sc_hd__dfrtp_4
X_15939_ _03402_ net350 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13852__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16439__X _02400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14895__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_305_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09460_ _03697_ _03700_ _03701_ _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_78_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18658_ clknet_leaf_60_clk _01075_ _00395_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[76\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16397__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17609_ net1914 _03020_ net429 vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15503__B _06573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09391_ net1135 net787 vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__or2_1
XANTENNA__18775__CLK clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_294_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18589_ clknet_leaf_31_clk _01009_ _00326_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[58\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_175_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_236_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09501__B game.CPU.applesa.ab.check_walls.above.walls\[52\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16149__A2 _01730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout134_A _02234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13958__B game.CPU.applesa.ab.check_walls.above.walls\[178\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11918__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19348__D game.CPU.applesa.twoapples.absxs.next_head\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18603__Q game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13383__A2 _07256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout301_A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16857__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_325_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09229__A game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11478__B net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09339__A1 net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19400__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09339__B2 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13974__A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_247_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_245_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1210_A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16350__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout101 net110 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1308_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout112 _02278_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_196_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout123 _02597_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_273_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15237__Y _08799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout134 _02234_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_261_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout145 net148 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout670_A _08799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14141__Y _08015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_X net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout156 net159 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_4
Xfanout167 net170 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_6
XANTENNA__16085__B2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A game.CPU.applesa.ab.apple_possible\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_226_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_346_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout189 net191 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_4
XANTENNA__19550__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ net1096 _03233_ _03965_ _03969_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__a211o_1
XANTENNA__13843__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16349__X _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17034__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09658_ net902 game.CPU.applesa.ab.check_walls.above.walls\[174\] game.CPU.applesa.ab.check_walls.above.walls\[175\]
+ net906 _03896_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_336_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09589_ net912 game.CPU.applesa.ab.check_walls.above.walls\[16\] net827 net908 vssd1
+ vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_258_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11620_ _05508_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11551_ game.CPU.applesa.ab.check_walls.above.walls\[195\] net762 vssd1 vssd1 vccd1
+ vccd1 _05440_ sky130_fd_sc_hd__xnor2_2
XANTENNA_clkbuf_leaf_69_clk_X clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_336_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16525__A net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_231_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13501__X _07375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10502_ game.CPU.applesa.ab.absxs.body_x\[79\] _04623_ _04624_ game.CPU.applesa.ab.absxs.body_x\[75\]
+ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__a22o_1
X_14270_ game.CPU.applesa.ab.absxs.body_y\[50\] net953 vssd1 vssd1 vccd1 vccd1 _08144_
+ sky130_fd_sc_hd__xnor2_1
X_11482_ net565 _05364_ _05368_ _05370_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__o211a_1
XANTENNA__16560__A2 _02481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20047__A game.CPU.applesa.ab.good_collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13221_ game.writer.tracker.frame\[388\] game.writer.tracker.frame\[389\] net1038
+ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__mux2_1
XANTENNA__13374__A2 _06710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10433_ game.CPU.bodymain1.Direction\[0\] _04573_ _04576_ vssd1 vssd1 vccd1 vccd1
+ _01220_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09578__B2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_268_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14045__A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_347_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11384__A2_N net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_249_Right_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13152_ net498 _07023_ _07025_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__a21o_1
XANTENNA__11388__B net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ game.CPU.walls.rand_wall.input2 game.CPU.walls.rand_wall.counter2\[0\] vssd1
+ vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__nor2_1
XFILLER_0_249_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19080__CLK net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12103_ _05989_ _05988_ _05987_ _05986_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_131_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_237_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17356__A _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13884__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13083_ game.writer.tracker.frame\[204\] game.writer.tracker.frame\[205\] net1010
+ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__mux2_1
X_17960_ net647 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__inv_2
XANTENNA__16260__A net248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10295_ net1450 _04473_ _04480_ game.CPU.applesa.ab.start_enable vssd1 vssd1 vccd1
+ vccd1 _01313_ sky130_fd_sc_hd__a22o_1
XFILLER_0_276_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18648__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08978__A game.CPU.applesa.ab.absxs.body_x\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16911_ _02322_ _02636_ net728 vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__o21a_1
X_12034_ game.CPU.applesa.ab.check_walls.above.walls\[140\] net551 vssd1 vssd1 vccd1
+ vccd1 _05921_ sky130_fd_sc_hd__or2_1
X_17891_ net620 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__inv_2
XANTENNA__13095__S net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19630_ clknet_leaf_27_clk game.writer.tracker.next_frame\[225\] net1309 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[225\] sky130_fd_sc_hd__dfrtp_1
X_16842_ game.writer.tracker.frame\[236\] _02616_ vssd1 vssd1 vccd1 vccd1 _02617_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_217_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_256_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout690 net691 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_205_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19561_ clknet_leaf_37_clk game.writer.tracker.next_frame\[156\] net1349 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[156\] sky130_fd_sc_hd__dfrtp_1
X_16773_ _02431_ net64 _02593_ net1960 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[190\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_109_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13985_ net985 game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1 vccd1
+ vccd1 _07859_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09502__A1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_358_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18512_ net580 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_358_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ net510 _06809_ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__or2_1
XFILLER_0_232_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_220_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15724_ game.CPU.applesa.ab.absxs.body_y\[55\] net435 vssd1 vssd1 vccd1 vccd1 _01736_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__09502__B2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19492_ clknet_leaf_24_clk game.writer.tracker.next_frame\[87\] net1338 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[87\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_272_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09602__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18443_ net592 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ game.writer.tracker.frame\[292\] game.writer.tracker.frame\[293\] net988
+ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__mux2_1
X_15655_ game.CPU.applesa.ab.check_walls.above.walls\[52\] net342 vssd1 vssd1 vccd1
+ vccd1 _01667_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14606_ _08460_ _08461_ net268 vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[6\]
+ sky130_fd_sc_hd__and3b_1
X_11818_ net750 _05322_ _05703_ _05705_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__a211oi_1
X_18374_ net598 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__inv_2
XANTENNA__15042__C net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15586_ game.CPU.applesa.ab.check_walls.above.walls\[32\] net271 vssd1 vssd1 vccd1
+ vccd1 _01598_ sky130_fd_sc_hd__nand2_1
XFILLER_0_334_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12798_ game.writer.tracker.frame\[342\] game.writer.tracker.frame\[343\] net1028
+ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_306_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17325_ net2002 net733 _02763_ _02428_ _02275_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[572\]
+ sky130_fd_sc_hd__a32o_1
X_14537_ _06547_ _06548_ _08410_ net556 vssd1 vssd1 vccd1 vccd1 game.writer.control.next\[0\]
+ sky130_fd_sc_hd__o2bb2a_1
X_11749_ game.CPU.applesa.ab.check_walls.above.walls\[174\] net300 net391 net785 vssd1
+ vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12963__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17256_ net135 net145 _02291_ net719 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__o31a_1
X_14468_ net1270 net859 net853 game.CPU.applesa.ab.absxs.body_y\[62\] vssd1 vssd1
+ vccd1 vccd1 _08342_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16551__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12682__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09569__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19423__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13419_ _06649_ _07002_ _07004_ _07003_ net504 net696 vssd1 vssd1 vccd1 vccd1 _07293_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09569__B2 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16207_ _01601_ _01602_ _01603_ _01608_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__or4_1
XANTENNA__12799__S1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17187_ _02492_ net77 _02727_ net1794 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[470\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_299_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_231_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14399_ game.CPU.applesa.ab.absxs.body_y\[69\] net962 vssd1 vssd1 vccd1 vccd1 _08273_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__16839__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12573__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13770__C1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_297_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16138_ _01664_ _02136_ _02140_ _02141_ _02149_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__o41a_1
XPHY_EDGE_ROW_216_Right_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15993__B net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_295_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13748__S0 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08960_ game.CPU.apple_location\[1\] vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__inv_2
X_16069_ game.CPU.applesa.ab.absxs.body_y\[87\] net431 vssd1 vssd1 vccd1 vccd1 _02081_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_5_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_255_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13522__C1 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10930__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14402__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17264__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19828_ clknet_leaf_38_clk game.writer.tracker.next_frame\[423\] net1333 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[423\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10887__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_320_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14078__B1 game.CPU.applesa.ab.YMAX\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19759_ clknet_leaf_26_clk game.writer.tracker.next_frame\[354\] net1313 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[354\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_242_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12697__X _06571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18097__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17016__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ _03751_ _03752_ _03753_ _03754_ _03750_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__a221o_1
XFILLER_0_223_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09443_ net1135 net791 vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11761__B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout251_A _05210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout349_A game.CPU.walls.rand_wall.abduyd.next_wall\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09374_ _03609_ _03611_ _03614_ _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__or4_1
XANTENNA__16790__A2 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14250__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13969__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1160_A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_331_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09885__C _04123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16064__B net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout304_X net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11367__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12564__B1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1046_X net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19916__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17098__A3 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09980__A1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14152__X _08026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16080__A game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1213_X net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10590__A2 _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_258_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10080_ _04286_ _04287_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_273_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_342_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14069__B1 _03380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12113__A game.CPU.applesa.ab.check_walls.above.walls\[53\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12619__A1 net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11952__A net569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ net514 _07639_ _07640_ _07643_ net216 vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__a311o_1
XFILLER_0_97_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10982_ _03267_ net413 vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_241_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12721_ _06572_ _06593_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15143__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11842__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15440_ _08921_ _08928_ _01466_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__o21ai_1
X_12652_ game.CPU.applesa.ab.absxs.body_x\[6\] net371 game.CPU.applesa.twoapples.absxs.next_head\[5\]
+ _03216_ _06451_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_318_Right_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_34_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14241__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_356_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16781__A2 _02454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16526__Y _02465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11055__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ game.CPU.applesa.ab.check_walls.above.walls\[97\] net771 vssd1 vssd1 vccd1
+ vccd1 _05492_ sky130_fd_sc_hd__xor2_1
XANTENNA__19446__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15371_ _08908_ _08912_ vssd1 vssd1 vccd1 vccd1 _08913_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_178_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ game.CPU.applesa.ab.absxs.body_x\[11\] net531 vssd1 vssd1 vccd1 vccd1 _06460_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__16255__A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_191_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17110_ net160 _02434_ net81 _02705_ net1565 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[415\]
+ sky130_fd_sc_hd__a32o_1
X_14322_ _08186_ _08187_ _08193_ _08195_ vssd1 vssd1 vccd1 vccd1 _08196_ sky130_fd_sc_hd__or4_1
X_18090_ net590 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__inv_2
X_11534_ _05420_ _05421_ _05422_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__or3_2
XFILLER_0_324_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16533__A2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_312_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17041_ _02396_ _02678_ _02683_ game.writer.tracker.frame\[368\] vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[368\] sky130_fd_sc_hd__a22o_1
XANTENNA__13347__A2 _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11399__A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14253_ game.CPU.applesa.ab.absxs.body_y\[23\] net941 vssd1 vssd1 vccd1 vccd1 _08127_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_351_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11465_ net777 _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13204_ game.writer.tracker.frame\[432\] game.writer.tracker.frame\[433\] net1035
+ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_170_Left_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19596__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ game.CPU.randy.f1.state\[0\] _04558_ _04557_ net931 vssd1 vssd1 vccd1 vccd1
+ _04562_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14184_ game.CPU.applesa.ab.absxs.body_y\[18\] net951 vssd1 vssd1 vccd1 vccd1 _08058_
+ sky130_fd_sc_hd__xor2_1
X_11396_ net778 _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16261__Y _02267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_267_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13135_ game.writer.tracker.frame\[164\] game.writer.tracker.frame\[165\] net1005
+ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__mux2_1
XANTENNA__09971__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10347_ _04487_ _04486_ game.CPU.randy.f1.a1.count\[0\] vssd1 vssd1 vccd1 vccd1 _01290_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__16836__A3 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18992_ net1197 _00218_ _00663_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_292_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_280_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_237_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13066_ game.writer.tracker.frame\[210\] game.writer.tracker.frame\[211\] net1026
+ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__mux2_1
X_17943_ net653 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__inv_2
X_10278_ _04391_ _04457_ _04462_ _04470_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__o211a_1
XANTENNA__19074__Q game.CPU.applesa.ab.check_walls.above.walls\[119\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12017_ game.CPU.applesa.ab.check_walls.above.walls\[44\] net554 vssd1 vssd1 vccd1
+ vccd1 _05904_ sky130_fd_sc_hd__nand2_1
X_17874_ net636 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__inv_2
XANTENNA__15037__C game.CPU.applesa.ab.check_walls.above.walls\[65\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17797__B2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_144_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19613_ clknet_leaf_20_clk game.writer.tracker.next_frame\[208\] net1310 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[208\] sky130_fd_sc_hd__dfrtp_1
X_16825_ _02362_ net143 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__and2b_1
XANTENNA__17261__A3 _02389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13807__B1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_232_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19544_ clknet_leaf_48_clk game.writer.tracker.next_frame\[139\] net1294 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[139\] sky130_fd_sc_hd__dfrtp_1
X_16756_ _02408_ net64 _02587_ net1744 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[179\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17549__A1 net1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13968_ _07837_ _07839_ _07841_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__or3_1
XANTENNA__12677__B net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_204_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15707_ game.CPU.applesa.ab.check_walls.above.walls\[152\] net269 vssd1 vssd1 vccd1
+ vccd1 _01719_ sky130_fd_sc_hd__or2_1
XFILLER_0_347_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12919_ net213 _06673_ net283 vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__a21o_1
X_19475_ clknet_leaf_19_clk game.writer.tracker.next_frame\[70\] net1335 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[70\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_278_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16687_ _02257_ _02280_ net98 net718 vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__o31a_1
X_13899_ net942 net816 vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_291_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_236_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18426_ net610 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__inv_2
X_15638_ game.CPU.applesa.ab.absxs.body_x\[81\] net471 vssd1 vssd1 vccd1 vccd1 _01650_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15988__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16772__A2 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16436__Y _02398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_302_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18357_ net596 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__inv_2
X_15569_ game.wr _01580_ _08877_ vssd1 vssd1 vccd1 vccd1 game.writer.updater.update.next\[2\]
+ sky130_fd_sc_hd__a21o_1
X_17308_ net1929 net723 _02759_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[559\]
+ sky130_fd_sc_hd__and3_1
X_09090_ game.CPU.applesa.ab.absxs.body_y\[57\] vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__inv_2
XANTENNA__18813__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19939__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18288_ net618 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16524__A2 _02462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17239_ _02549_ net79 _02740_ net1885 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[509\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_303_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16315__D net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18380__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_330_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_302_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15509__A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16827__A3 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09992_ game.CPU.apple_location\[7\] net1458 _04207_ vssd1 vssd1 vccd1 vccd1 _01372_
+ sky130_fd_sc_hd__mux2_1
X_08943_ net1089 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_244_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout299_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__A1 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__B2 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_327_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_243_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19319__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1006_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17252__A3 _02280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13971__B game.CPU.applesa.ab.check_walls.above.walls\[82\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15799__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout466_A net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16460__B2 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12587__B net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16059__B net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11491__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19469__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17004__A3 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout254_X net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ net1147 net798 vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__or2_1
XFILLER_0_338_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_255_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15898__B net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16763__A2 _02331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11037__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09357_ net1098 _03484_ _03487_ net1128 _03599_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14147__X _08021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09288_ net1137 net809 vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_97_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16515__A2 _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17712__A1 net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10260__A1 game.CPU.applesa.ab.XMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10260__B2 game.CPU.applesa.ab.XMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18290__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12108__A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ _04991_ _04992_ _05138_ _05139_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09402__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17618__B net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_344_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout888_X net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ net1168 net765 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11181_ game.CPU.applesa.ab.absxs.body_x\[78\] net410 vssd1 vssd1 vccd1 vccd1 _05071_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__14323__A game.CPU.applesa.ab.absxs.body_x\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_274_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09417__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ game.CPU.randy.f1.c1.count\[3\] game.CPU.randy.f1.c1.count\[4\] vssd1 vssd1
+ vccd1 vccd1 _04327_ sky130_fd_sc_hd__nand2_1
XANTENNA__15138__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14042__B net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17228__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09705__B2 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ _04225_ _04270_ _04228_ _04217_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__o211a_1
X_14940_ _08715_ _08716_ vssd1 vssd1 vccd1 vccd1 _08717_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_237_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14871_ net1433 _08655_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[18\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_214_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16610_ net202 _02453_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__nor2_4
XFILLER_0_202_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15154__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11682__A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13822_ net216 _07691_ net280 vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_106_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17590_ game.CPU.kyle.L1.cnt_20ms\[1\] game.CPU.kyle.L1.cnt_20ms\[0\] vssd1 vssd1
+ vccd1 vccd1 _03010_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12497__B net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_355_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16541_ net113 _02473_ net716 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__o21a_1
X_13753_ _07623_ _07626_ net204 vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__mux2_1
XANTENNA__11276__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10965_ game.CPU.applesa.ab.absxs.body_y\[117\] net542 vssd1 vssd1 vccd1 vccd1 _04855_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10298__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12704_ _06569_ _06577_ _06568_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__a21oi_2
X_19260_ clknet_leaf_57_clk _01328_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.count_luck\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_13684_ _07556_ _07557_ net487 vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__mux2_1
X_16472_ net167 net195 _02297_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__and3_4
XANTENNA__08991__A game.CPU.applesa.ab.absxs.body_x\[55\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10896_ game.CPU.applesa.ab.check_walls.collision_up _04797_ vssd1 vssd1 vccd1 vccd1
+ _04798_ sky130_fd_sc_hd__or2_1
XANTENNA__14214__B1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18211_ net666 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__inv_2
X_15423_ game.writer.updater.commands.cmd_num\[1\] _01436_ game.writer.updater.commands.cmd_num\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12635_ _06508_ _06509_ _06510_ _06511_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__or4_1
X_19191_ clknet_leaf_46_clk net348 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.x_final\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__15601__B net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15354_ game.writer.updater.commands.count\[6\] game.writer.updater.commands.count\[5\]
+ _08895_ game.writer.updater.commands.count\[7\] vssd1 vssd1 vccd1 vccd1 _08896_
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18142_ net631 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__inv_2
X_12566_ _03286_ game.CPU.applesa.twoapples.absxs.next_head\[2\] net361 game.CPU.applesa.ab.absxs.body_y\[116\]
+ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_297_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire140 _02569_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_1
XANTENNA__18986__CLK net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14305_ game.CPU.applesa.ab.absxs.body_x\[28\] net1070 vssd1 vssd1 vccd1 vccd1 _08179_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_108_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11517_ net832 _05210_ _05396_ net193 vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18073_ net658 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__inv_2
X_15285_ _08817_ _08832_ vssd1 vssd1 vccd1 vccd1 _08837_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12497_ game.CPU.applesa.ab.absxs.body_x\[65\] net379 vssd1 vssd1 vccd1 vccd1 _06374_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12528__B1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13725__C1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold209 game.writer.tracker.frame\[427\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
X_17024_ net1466 _02677_ _02679_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[355\]
+ sky130_fd_sc_hd__a21o_1
X_14236_ game.CPU.applesa.ab.absxs.body_x\[113\] net1067 vssd1 vssd1 vccd1 vccd1 _08110_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11448_ net779 _05336_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__xor2_1
XFILLER_0_278_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_308_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11200__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18701__Q game.CPU.applesa.ab.absxs.body_x\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16809__A3 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14167_ game.CPU.applesa.ab.absxs.body_y\[104\] net989 vssd1 vssd1 vccd1 vccd1 _08041_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_150_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_237_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14233__A game.CPU.applesa.ab.absxs.body_x\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11379_ game.CPU.applesa.ab.check_walls.above.walls\[177\] net770 vssd1 vssd1 vccd1
+ vccd1 _05268_ sky130_fd_sc_hd__xnor2_1
X_13118_ net696 _06991_ _06988_ net204 vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__o211a_1
XANTENNA__11576__B net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14098_ _07970_ _07971_ _07964_ _07969_ vssd1 vssd1 vccd1 vccd1 _07972_ sky130_fd_sc_hd__a211o_1
XANTENNA__15048__B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18975_ net1198 _00200_ _00646_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_294_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16690__A1 _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13049_ game.writer.tracker.frame\[252\] game.writer.tracker.frame\[253\] net1031
+ vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17926_ net606 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__inv_2
XFILLER_0_294_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1260 game.CPU.randy.f1.state\[5\] vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__clkbuf_2
Xfanout1271 net1273 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__buf_4
XANTENNA__17234__A3 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17857_ game.writer.updater.commands.count\[12\] game.writer.updater.commands.count\[11\]
+ _03172_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__and3_1
Xfanout1282 net1283 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12688__A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13283__S net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_280_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1293 net1360 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__buf_2
XFILLER_0_353_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19611__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16442__A1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11592__A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15064__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16808_ _02494_ net99 net727 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__o21a_1
Xclkbuf_3_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__14453__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17788_ net757 game.CPU.applesa.twomode.counter_flip vssd1 vssd1 vccd1 vccd1 _01385_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__16993__A2 net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10479__Y _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09062__A game.CPU.applesa.ab.absxs.body_y\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19527_ clknet_leaf_22_clk game.writer.tracker.next_frame\[122\] net1342 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[122\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16739_ _02370_ _02561_ net719 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__o21a_1
XANTENNA__12200__B net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_313_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_347_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19458_ clknet_leaf_39_clk game.writer.tracker.next_frame\[53\] net1352 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[53\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14205__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19761__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09880__B1 _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16607__B _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09211_ game.CPU.applesa.ab.check_walls.above.walls\[155\] vssd1 vssd1 vccd1 vccd1
+ _03460_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13559__A2 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18409_ net602 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__inv_2
XANTENNA__10447__D_N net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19389_ clknet_leaf_4_clk _01395_ _00969_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.snake_head_x\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_146_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09142_ game.CPU.applesa.ab.check_walls.above.walls\[25\] vssd1 vssd1 vccd1 vccd1
+ _03391_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_288_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09073_ game.CPU.applesa.ab.absxs.body_y\[114\] vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15705__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_315_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17170__A2 _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_287_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout214_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16623__A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_250_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13716__C1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_330_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13458__S net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19356__D game.CPU.applesa.twoapples.absxs.next_head\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13731__A2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12215__X _06101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10671__A _04594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11742__A1 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19141__CLK net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09975_ net1261 _04201_ _04202_ _04158_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__o211a_1
XANTENNA__18709__CLK clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13982__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_243_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_164_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1009_X net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout750_A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19291__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18859__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16984__A2 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13798__A2 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13342__S1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1280_X net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10750_ game.CPU.applesa.ab.absxs.body_y\[113\] _04663_ _04664_ game.CPU.applesa.ab.absxs.body_y\[109\]
+ vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__a22o_1
XANTENNA__15702__A game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_338_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_326_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16736__A2 _02524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12470__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_338_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09409_ net1097 game.CPU.applesa.ab.check_walls.above.walls\[129\] vssd1 vssd1 vccd1
+ vccd1 _03652_ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10681_ game.CPU.applesa.ab.absxs.body_x\[11\] _04689_ _04707_ game.CPU.applesa.ab.absxs.body_x\[7\]
+ vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_326_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12420_ game.CPU.applesa.ab.absxs.body_y\[33\] net523 net363 game.CPU.applesa.ab.absxs.body_y\[32\]
+ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_350_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_341_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_303_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12351_ game.CPU.applesa.ab.absxs.body_y\[76\] net360 vssd1 vssd1 vccd1 vccd1 _06228_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_306_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17161__A2 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12037__A1_N net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13707__C1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10784__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11302_ _04973_ _05146_ _05162_ _05191_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.collision
+ sky130_fd_sc_hd__nand4_4
X_15070_ net1216 net1238 game.CPU.applesa.ab.check_walls.above.walls\[98\] vssd1 vssd1
+ vccd1 vccd1 _00095_ sky130_fd_sc_hd__and3_1
X_12282_ game.CPU.applesa.ab.check_walls.above.walls\[133\] net547 vssd1 vssd1 vccd1
+ vccd1 _06168_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14021_ _07885_ _07889_ _07892_ _07894_ vssd1 vssd1 vccd1 vccd1 _07895_ sky130_fd_sc_hd__or4_2
X_11233_ game.CPU.applesa.ab.absxs.body_x\[15\] net545 vssd1 vssd1 vccd1 vccd1 _05123_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__15149__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13722__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10581__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12125__X _06012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11733__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10536__A2 _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_264_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09147__A game.CPU.applesa.ab.check_walls.above.walls\[32\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16121__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ game.CPU.applesa.ab.absxs.body_y\[50\] net539 _04819_ game.CPU.applesa.ab.absxs.body_y\[48\]
+ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__a22o_1
XANTENNA__14988__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19634__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16672__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10115_ _04317_ net1475 _04311_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_186_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18760_ clknet_leaf_12_clk _01177_ _00497_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[54\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13486__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11095_ _03339_ net404 vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__xnor2_1
X_15972_ game.CPU.applesa.ab.absxs.body_x\[64\] net271 vssd1 vssd1 vccd1 vccd1 _01984_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__08986__A game.CPU.applesa.ab.absxs.body_x\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09434__X _03677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17711_ _04255_ _04471_ net1166 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_303_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14923_ _08657_ _08677_ _08699_ vssd1 vssd1 vccd1 vccd1 _08700_ sky130_fd_sc_hd__or3b_1
X_10046_ net846 vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__inv_2
X_18691_ clknet_leaf_65_clk _01108_ _00428_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[33\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_262_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold70 game.CPU.applesa.ab.count\[3\] vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14500__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold81 game.writer.tracker.frame\[355\] vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_203_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17642_ game.CPU.kyle.L1.cnt_500hz\[4\] _08802_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__or2_1
Xhold92 net46 vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_264_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14854_ game.CPU.randy.f1.c1.count\[11\] game.CPU.randy.f1.c1.count\[10\] _08645_
+ vssd1 vssd1 vccd1 vccd1 _08647_ sky130_fd_sc_hd__and3_1
XANTENNA__14435__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19784__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16975__A2 _02452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_199_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13805_ net513 _07675_ _07676_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__and3_1
XFILLER_0_202_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17573_ _02844_ _02870_ _02875_ _02996_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__or4_1
X_14785_ _03512_ _08603_ vssd1 vssd1 vccd1 vccd1 _08604_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11997_ net825 net297 net291 game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1
+ vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__a22o_1
XANTENNA__16708__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_230_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19312_ net1163 _00036_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.out_random_2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16524_ net125 _02462_ net558 vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_275_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15612__A game.CPU.applesa.ab.absxs.body_x\[35\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13736_ net212 _07603_ net283 vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__o21a_1
XFILLER_0_202_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10948_ _03247_ net408 vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16727__A2 _02434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_280_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_217_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09610__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19243_ clknet_leaf_17_clk _00074_ _00881_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__19014__CLK net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_329_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16455_ net185 net118 _02412_ _02406_ net1888 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[53\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__15935__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13667_ net245 _07539_ _07524_ net183 vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__o211a_1
X_10879_ game.CPU.applesa.ab.apple_possible\[7\] _04780_ vssd1 vssd1 vccd1 vccd1 _04781_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15406_ game.writer.updater.commands.cmd_num\[3\] _08935_ _01433_ _08911_ vssd1 vssd1
+ vccd1 vccd1 _01434_ sky130_fd_sc_hd__a22o_1
XFILLER_0_213_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19174_ clknet_leaf_4_clk _01293_ _00836_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12618_ _03235_ game.CPU.applesa.twoapples.absxs.next_head\[3\] game.CPU.applesa.twoapples.absxs.next_head\[6\]
+ _03300_ _06231_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_314_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16386_ net244 net236 _02296_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__or3_4
X_13598_ game.writer.tracker.frame\[297\] game.writer.tracker.frame\[299\] game.writer.tracker.frame\[300\]
+ game.writer.tracker.frame\[298\] net973 net988 vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__mux4_1
XANTENNA__12844__S0 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18125_ net577 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__inv_2
X_15337_ _06546_ _08878_ vssd1 vssd1 vccd1 vccd1 _08879_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12549_ _03250_ net376 vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_269_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10775__A2 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19164__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11972__B2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18056_ net653 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__inv_2
XANTENNA_1 _02179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ _08823_ vssd1 vssd1 vccd1 vccd1 _08824_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17007_ _02497_ net84 _02673_ net1804 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[344\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14910__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15059__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14219_ game.CPU.applesa.ab.absxs.body_y\[40\] net869 net860 game.CPU.applesa.ab.absxs.body_y\[43\]
+ vssd1 vssd1 vccd1 vccd1 _08093_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_286_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14910__B2 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15199_ _03524_ game.CPU.applesa.normal1.number\[0\] game.CPU.applesa.normal1.number\[1\]
+ vssd1 vssd1 vccd1 vccd1 _08768_ sky130_fd_sc_hd__or3_1
XANTENNA__16730__X _02579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__A2 _04609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_300_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout508 net515 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_228_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14898__A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout519 net522 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__buf_4
XFILLER_0_308_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09760_ net923 game.CPU.applesa.ab.check_walls.above.walls\[26\] game.CPU.applesa.ab.check_walls.above.walls\[29\]
+ net899 vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a22o_1
XANTENNA__12910__S net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18958_ net1200 _00221_ _00629_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_17909_ net668 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__inv_2
X_09691_ net1109 game.CPU.applesa.ab.absxs.body_x\[4\] vssd1 vssd1 vccd1 vccd1 _03934_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__13572__S1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18889_ clknet_leaf_1_clk _01261_ vssd1 vssd1 vccd1 vccd1 game.CPU.kyle.L1.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xfanout1090 net1091 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__buf_4
XANTENNA__16415__B2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17612__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16122__A2_N net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_317_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13324__S1 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout164_A net165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_239_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_335_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_252_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout429_A _00293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19507__CLK clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_335_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ net990 vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13977__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17143__A2 _02415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout217_X net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1240_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10766__A2 _04673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11963__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ game.CPU.applesa.ab.absxs.body_y\[62\] vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_328_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19437__Q game.writer.tracker.frame\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_288_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16072__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19657__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold540 game.writer.tracker.frame\[229\] vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 game.writer.tracker.frame\[540\] vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11715__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1126_X net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 game.writer.tracker.frame\[14\] vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10832__C _04737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold573 game.writer.tracker.frame\[456\] vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 game.writer.tracker.frame\[338\] vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_275_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold595 game.CPU.clock1.counter\[16\] vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_291_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout965_A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11191__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12820__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_290_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09958_ net1146 _04186_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__or2_1
XANTENNA__18681__CLK clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11944__B net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ _03999_ _04005_ _04131_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__o21a_2
XANTENNA__16406__B2 _01516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11920_ _05800_ _05804_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__or3_1
XANTENNA__12121__A game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_339_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12419__A2_N net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11851_ net570 _05364_ _05368_ _05369_ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__17631__B net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout920_X net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16830__A_N net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_352_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12979__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14974__C game.CPU.applesa.ab.check_walls.above.walls\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10802_ game.CPU.applesa.ab.absxs.body_y\[27\] _04695_ _04698_ game.CPU.applesa.ab.absxs.body_y\[23\]
+ vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__a22o_1
XANTENNA__11960__A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14570_ _04482_ _08432_ _08433_ game.CPU.clock1.game_state\[0\] vssd1 vssd1 vccd1
+ vccd1 game.CPU.state1.Qn\[0\] sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_123_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ game.CPU.applesa.ab.check_walls.above.walls\[84\] net392 net301 net809 _05667_
+ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__o221a_1
XFILLER_0_184_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13521_ net279 _07345_ _07349_ net241 vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__o31a_1
XFILLER_0_177_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15151__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ game.CPU.applesa.ab.absxs.body_y\[22\] _04645_ _04652_ game.CPU.applesa.ab.absxs.body_y\[18\]
+ vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__a22o_1
XANTENNA__14048__A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19187__CLK net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13452_ net214 _07321_ _07325_ net285 vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__o211a_1
X_16240_ _06573_ _02245_ _02247_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_192_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14196__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10664_ _04174_ _04583_ _04606_ net848 vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a31o_4
XFILLER_0_165_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_341_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12403_ game.CPU.applesa.ab.absxs.body_x\[52\] net382 vssd1 vssd1 vccd1 vccd1 _06280_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_341_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13887__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13383_ _07209_ _07256_ _07255_ net177 vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__o211a_1
X_16171_ _03275_ net347 net432 game.CPU.applesa.ab.absxs.body_y\[35\] _02124_ vssd1
+ vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a221o_1
X_10595_ _03229_ net263 vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__nor2_1
XANTENNA__17134__A2 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12334_ game.CPU.applesa.twoapples.logic_enable _04237_ _06211_ vssd1 vssd1 vccd1
+ vccd1 _06214_ sky130_fd_sc_hd__a21o_2
X_15122_ net1208 net1233 game.CPU.applesa.ab.check_walls.above.walls\[150\] vssd1
+ vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_188_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13098__S net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19930_ clknet_leaf_33_clk game.writer.tracker.next_frame\[525\] net1302 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[525\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16893__A1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15053_ net1217 net1245 game.CPU.applesa.ab.check_walls.above.walls\[81\] vssd1 vssd1
+ vccd1 vccd1 _00275_ sky130_fd_sc_hd__and3_1
X_12265_ game.CPU.applesa.ab.check_walls.above.walls\[109\] net548 vssd1 vssd1 vccd1
+ vccd1 _06151_ sky130_fd_sc_hd__or2_1
XFILLER_0_160_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10509__A2 _04625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11706__A1 game.CPU.applesa.ab.check_walls.above.walls\[165\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14004_ net867 game.CPU.applesa.ab.check_walls.above.walls\[140\] game.CPU.applesa.ab.check_walls.above.walls\[136\]
+ net886 vssd1 vssd1 vccd1 vccd1 _07878_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_39_Left_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11216_ game.CPU.applesa.ab.absxs.body_x\[38\] net320 vssd1 vssd1 vccd1 vccd1 _05106_
+ sky130_fd_sc_hd__nand2_1
X_19861_ clknet_leaf_20_clk game.writer.tracker.next_frame\[456\] net1315 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[456\] sky130_fd_sc_hd__dfrtp_1
X_12196_ net825 net424 vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__xnor2_1
X_18812_ clknet_leaf_72_clk game.CPU.clock1.next_counter\[15\] _00549_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16645__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11147_ game.CPU.applesa.ab.absxs.body_x\[97\] net414 net411 game.CPU.applesa.ab.absxs.body_x\[98\]
+ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__a22o_1
XANTENNA__15607__A game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19792_ clknet_leaf_35_clk game.writer.tracker.next_frame\[387\] net1348 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[387\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13459__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12730__S net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09605__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18743_ clknet_leaf_10_clk _01160_ _00480_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_15955_ _03394_ net338 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__xnor2_1
X_11078_ game.CPU.applesa.ab.absxs.body_y\[43\] net397 vssd1 vssd1 vccd1 vccd1 _04968_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__19082__Q game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12131__A1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12131__B2 game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10029_ net1163 game.CPU.applesa.out_random_2\[6\] vssd1 vssd1 vccd1 vccd1 _04237_
+ sky130_fd_sc_hd__nand2_2
X_14906_ _08681_ _08682_ vssd1 vssd1 vccd1 vccd1 _08683_ sky130_fd_sc_hd__and2b_1
X_18674_ clknet_leaf_8_clk _01091_ _00411_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_223_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15886_ game.CPU.applesa.ab.check_walls.above.walls\[141\] net444 vssd1 vssd1 vccd1
+ vccd1 _01898_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15045__C game.CPU.applesa.ab.check_walls.above.walls\[73\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14408__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16948__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17070__A1 _02444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17625_ game.CPU.kyle.L1.cnt_20ms\[14\] game.CPU.kyle.L1.cnt_20ms\[13\] _03028_ vssd1
+ vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__and3_1
X_14837_ game.CPU.randy.f1.c1.count\[4\] _08635_ vssd1 vssd1 vccd1 vccd1 _08637_ sky130_fd_sc_hd__or2_1
XFILLER_0_175_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17556_ _02778_ net427 _02840_ _02937_ _02981_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__a32o_1
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14768_ game.CPU.randy.counter1.count\[7\] game.CPU.randy.counter1.count\[5\] net266
+ vssd1 vssd1 vccd1 vccd1 _08589_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12434__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16507_ net1769 _02446_ _02450_ net128 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[66\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_317_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13719_ _07591_ _07592_ net478 vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__mux2_1
X_17487_ _02883_ _02915_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14699_ _08505_ _08516_ _08524_ _08515_ vssd1 vssd1 vccd1 vccd1 _08538_ sky130_fd_sc_hd__or4b_1
XFILLER_0_316_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19226_ net1167 _01320_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.normal1.counter_normal
+ sky130_fd_sc_hd__dfxtp_1
X_16438_ _02247_ net237 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__or2_1
XANTENNA__14187__A2 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_288_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18554__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_310_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19157_ clknet_leaf_3_clk _01278_ _00828_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.counter2\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13934__A2 game.CPU.applesa.ab.check_walls.above.walls\[32\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12905__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16369_ _06573_ _02231_ _02313_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__or3b_2
XANTENNA__17125__A2 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10748__A2 _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18108_ net628 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__inv_2
X_19088_ net1177 _00125_ _00759_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[133\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10933__B net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18039_ net602 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__inv_2
XANTENNA__12206__A game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout305 net307 vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_273_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16620__B net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout316 net318 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_2
XFILLER_0_319_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20001_ clknet_leaf_44_clk _01425_ net1300 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[16\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__buf_2
X_09812_ net1155 game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1 _04055_
+ sky130_fd_sc_hd__or2_1
Xfanout338 net339 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_2
XFILLER_0_272_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout349 game.CPU.walls.rand_wall.abduyd.next_wall\[2\] vssd1 vssd1 vccd1 vccd1
+ net349 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_323_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09743_ net1141 game.CPU.applesa.ab.check_walls.above.walls\[70\] vssd1 vssd1 vccd1
+ vccd1 _03986_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_161_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout281_A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout379_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_198_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09674_ net1085 net1265 vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__nand2_1
XFILLER_0_335_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13870__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17061__A1 _02435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13870__B2 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10684__A1 game.CPU.applesa.ab.absxs.body_x\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16348__A net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1190_A game.CPU.walls.rand_wall.good_spot vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout167_X net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_327_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16067__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16635__X _02535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_308_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_172_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_308_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_350_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_323_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout501_X net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17116__A2 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12815__S net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_X net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10739__A2 _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ game.CPU.applesa.ab.absxs.body_y\[8\] vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__inv_2
XFILLER_0_350_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10380_ net1144 _03205_ _03206_ net1096 _04532_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14315__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14003__A1_N net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09039_ game.CPU.applesa.ab.absxs.body_x\[116\] vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__inv_2
XANTENNA__17907__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13689__A1 _07554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13689__B2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12050_ net817 net553 vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__or2_1
Xhold370 game.writer.tracker.frame\[76\] vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14350__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold381 game.writer.tracker.frame\[284\] vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17626__B net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold392 game.writer.tracker.frame\[199\] vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16530__B _02340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_261_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout968_X net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16627__A1 _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11164__A2 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ _03242_ net406 net402 _03309_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_183_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout850 _04157_ vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09425__A net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout861 net863 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_4
XANTENNA__11674__B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout872 _03374_ vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_4
XANTENNA__15146__B net1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout883 net884 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_125_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout894 net895 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_300_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16029__A2_N net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15740_ game.CPU.applesa.ab.check_walls.above.walls\[173\] net444 vssd1 vssd1 vccd1
+ vccd1 _01752_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_245_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12952_ net481 _06825_ _06824_ net224 vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__o211a_1
XANTENNA__13861__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14985__B net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17052__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17052__B2 game.writer.tracker.frame\[376\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10675__A1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ game.CPU.applesa.ab.check_walls.above.walls\[44\] net394 _05782_ _05783_
+ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__o2111a_1
X_15671_ _03437_ net343 vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__nor2_1
X_12883_ game.writer.tracker.frame\[16\] game.writer.tracker.frame\[17\] net1006 vssd1
+ vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17410_ game.CPU.speed1.Qa\[0\] game.CPU.speed1.Qa\[2\] vssd1 vssd1 vccd1 vccd1 _02840_
+ sky130_fd_sc_hd__or2_2
XANTENNA__15162__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11690__A net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_261_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14622_ _08470_ _08471_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[12\]
+ sky130_fd_sc_hd__nor2_1
X_18390_ net600 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
X_11834_ game.CPU.applesa.ab.check_walls.above.walls\[151\] net310 vssd1 vssd1 vccd1
+ vccd1 _05722_ sky130_fd_sc_hd__nand2_1
XANTENNA__13613__A1 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09160__A game.CPU.applesa.ab.check_walls.above.walls\[53\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_272_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18577__CLK clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17341_ _08751_ _08753_ _02769_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__a21o_1
X_14553_ game.CPU.walls.rand_wall.logic_enable _04253_ net1272 vssd1 vssd1 vccd1 vccd1
+ _08422_ sky130_fd_sc_hd__a21oi_1
X_11765_ _05269_ _05270_ _05651_ _05652_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__and4b_1
XANTENNA__19822__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13504_ net279 _07333_ _07334_ net241 vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__a31o_1
X_10716_ game.CPU.applesa.ab.absxs.body_y\[54\] _04609_ _04637_ game.CPU.applesa.ab.absxs.body_y\[50\]
+ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__a22o_1
X_17272_ net136 net70 _02328_ net733 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_194_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ net774 _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14484_ _08262_ _08267_ _08357_ _08141_ vssd1 vssd1 vccd1 vccd1 _08358_ sky130_fd_sc_hd__o211a_1
XFILLER_0_342_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13377__B1 _07250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19011_ net1202 _00239_ _00682_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[56\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16223_ net1693 _02232_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[1\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_136_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13435_ _06936_ _06967_ net686 vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__mux2_1
X_10647_ _04692_ game.CPU.applesa.ab.absxs.body_x\[42\] _04690_ vssd1 vssd1 vccd1
+ vccd1 _01113_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_311_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17107__A2 _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_299_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11927__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13366_ net213 _07235_ net283 vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__a21o_1
X_16154_ _01713_ _01714_ _01718_ _01719_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a22o_1
XANTENNA__19972__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10578_ _03255_ net234 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_47_Left_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14225__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15105_ net1204 net1231 net792 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12317_ _06080_ _06081_ _06082_ _06107_ _06202_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__o311a_1
X_13297_ net499 _07170_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__or2_1
XFILLER_0_239_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16085_ game.CPU.applesa.ab.check_walls.above.walls\[145\] net471 net430 net789 _02096_
+ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__o221a_1
XANTENNA__16721__A _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12026__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19913_ clknet_leaf_22_clk game.writer.tracker.next_frame\[508\] net1339 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[508\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_294_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12248_ net797 net418 vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__xnor2_1
X_15036_ net1219 net1244 game.CPU.applesa.ab.check_walls.above.walls\[64\] vssd1 vssd1
+ vccd1 vccd1 _00257_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_283_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_239_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14341__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16440__B _02400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19202__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16618__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_225_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11865__A game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_19844_ clknet_leaf_36_clk game.writer.tracker.next_frame\[439\] net1357 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[439\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_299_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12179_ _06039_ _06040_ _06041_ _06049_ _06065_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__o311a_1
XFILLER_0_286_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_247_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17291__A1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12483__A1_N game.CPU.applesa.ab.absxs.body_y\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09335__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19775_ clknet_leaf_26_clk game.writer.tracker.next_frame\[370\] net1312 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[370\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15056__B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16987_ net145 _02467_ net88 _02667_ net1472 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[330\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_266_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18726_ clknet_leaf_13_clk _01143_ _00463_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[108\]
+ sky130_fd_sc_hd__dfrtp_4
X_15938_ _01943_ _01945_ _01946_ _01949_ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17043__A1 _02398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_56_Left_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_250_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10666__A1 game.CPU.applesa.ab.absxs.body_x\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_305_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18657_ clknet_leaf_51_clk _01074_ _00394_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[71\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10666__B2 game.CPU.applesa.ab.absxs.body_x\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15869_ game.CPU.applesa.ab.absxs.body_y\[27\] net432 vssd1 vssd1 vccd1 vccd1 _01881_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17608_ game.CPU.kyle.L1.cnt_20ms\[8\] _03020_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__and2_1
XANTENNA__15072__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_175_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09390_ net1135 net787 vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_171_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_294_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18588_ clknet_leaf_31_clk _01008_ _00325_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[57\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12407__A2 game.CPU.applesa.twoapples.absxs.next_head\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17539_ net1243 _02845_ _02920_ _02964_ _02965_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__a2111o_1
XANTENNA__12983__X _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_236_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18383__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_321_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_352_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11105__A game.CPU.applesa.ab.absxs.body_x\[35\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__16554__B1 _02483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19209_ net1167 _00021_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_possible\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_6_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_332_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10944__A game.CPU.applesa.ab.absxs.body_x\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout127_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11918__B2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12040__B1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16857__A1 net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_325_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1036_A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16350__B net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_247_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13466__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout102 net103 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13540__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout113 net114 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__buf_4
Xfanout124 net129 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_4
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_4
XFILLER_0_196_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout146 net147 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
Xfanout157 net158 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17282__A1 net176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09245__A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16085__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout168 net170 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11494__B net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_260_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout663_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09726_ net891 game.CPU.applesa.ab.absxs.body_y\[84\] _03967_ _03968_ vssd1 vssd1
+ vccd1 vccd1 _03969_ sky130_fd_sc_hd__a211o_1
XFILLER_0_179_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10657__A1 game.CPU.applesa.ab.absxs.body_x\[33\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_96_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ net1089 game.CPU.applesa.ab.check_walls.above.walls\[170\] vssd1 vssd1 vccd1
+ vccd1 _03900_ sky130_fd_sc_hd__xor2_1
XANTENNA__11854__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_336_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19845__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09588_ net1112 _03386_ game.CPU.applesa.ab.check_walls.above.walls\[20\] net894
+ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_355_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_258_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1360_X net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_231_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11550_ _05436_ _05437_ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__or3_1
XANTENNA__19995__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16525__B _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Left_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10501_ net1080 _04623_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__nor2_2
XFILLER_0_162_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11481_ _04450_ _05365_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11909__A1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14326__A game.CPU.applesa.ab.absxs.body_y\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_323_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ net704 _07093_ _07090_ net230 vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__o211a_1
XFILLER_0_323_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_311_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10432_ _04563_ _04569_ _04573_ _04574_ game.CPU.bodymain1.main.pause_clk vssd1 vssd1
+ vccd1 vccd1 _04576_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_323_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12031__B1 _05894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11385__A2 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_347_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13151_ net514 _07024_ net689 vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__a21o_1
XFILLER_0_289_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10363_ game.CPU.walls.rand_wall.counter2\[4\] game.CPU.walls.rand_wall.counter2\[3\]
+ game.CPU.walls.rand_wall.counter2\[2\] _04524_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__or4_1
XFILLER_0_150_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12102_ _05301_ _05302_ _05304_ _05306_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__or4b_1
X_13082_ game.writer.tracker.frame\[208\] game.writer.tracker.frame\[209\] net1010
+ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__mux2_1
XANTENNA__15520__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10294_ _03494_ game.CPU.applesa.ab.x_final\[1\] game.CPU.applesa.ab.good_spot_next
+ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__and3_1
XFILLER_0_237_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13531__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16910_ _02486_ net95 _02645_ net1708 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[275\]
+ sky130_fd_sc_hd__a22o_1
X_12033_ game.CPU.applesa.ab.check_walls.above.walls\[140\] net551 vssd1 vssd1 vccd1
+ vccd1 _05920_ sky130_fd_sc_hd__nand2_1
XANTENNA__11685__A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_256_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15157__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_236_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17890_ net620 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__inv_2
XANTENNA__12133__X _06020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19375__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17273__A1 _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Left_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16841_ net131 _02299_ net142 _02616_ net1663 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[235\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_8_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14087__A1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14996__A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 net681 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14087__B2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout691 net692 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__buf_2
X_19560_ clknet_leaf_37_clk game.writer.tracker.next_frame\[155\] net1349 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[155\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12098__B1 _05977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16772_ _02429_ net64 _02593_ net1942 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[189\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13984_ _07854_ _07855_ _07856_ _07857_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__a22o_1
XANTENNA__17025__A1 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18511_ net580 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__inv_2
X_15723_ game.CPU.applesa.ab.absxs.body_y\[52\] net341 vssd1 vssd1 vccd1 vccd1 _01735_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__09502__A2 game.CPU.applesa.ab.check_walls.above.walls\[49\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_358_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12935_ _06719_ _06722_ net686 vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__mux2_1
X_19491_ clknet_leaf_23_clk game.writer.tracker.next_frame\[86\] net1339 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[86\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11845__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_358_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17576__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13405__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ net592 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__inv_2
XFILLER_0_272_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15654_ game.CPU.applesa.ab.check_walls.above.walls\[164\] net450 net472 game.CPU.applesa.ab.check_walls.above.walls\[161\]
+ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09602__B game.CPU.applesa.ab.absxs.body_x\[73\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_157_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12866_ game.writer.tracker.frame\[296\] game.writer.tracker.frame\[297\] net988
+ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14605_ game.CPU.clock1.counter\[5\] _08458_ game.CPU.clock1.counter\[6\] vssd1 vssd1
+ vccd1 vccd1 _08461_ sky130_fd_sc_hd__a21o_1
X_18373_ net598 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__inv_2
X_11817_ _05324_ _05704_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16275__X _02280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15585_ _01591_ _01594_ _01595_ _01596_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__or4_2
X_12797_ game.writer.tracker.frame\[338\] game.writer.tracker.frame\[339\] net1028
+ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17324_ net1905 net732 _02763_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[571\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__15620__A game.CPU.applesa.ab.check_walls.above.walls\[87\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14536_ _08406_ _08407_ _08409_ vssd1 vssd1 vccd1 vccd1 _08410_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_185_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_327_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11748_ _05619_ _05623_ _05625_ _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16000__A2 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17255_ net111 _02466_ _02744_ net1964 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[521\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10820__A1 game.CPU.applesa.ab.absxs.body_y\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14467_ _03239_ net1066 net859 net1270 vssd1 vssd1 vccd1 vccd1 _08341_ sky130_fd_sc_hd__o22a_1
XANTENNA__10820__B2 game.CPU.applesa.ab.absxs.body_y\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11679_ game.CPU.applesa.ab.check_walls.above.walls\[58\] game.CPU.applesa.ab.apple_possible\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__xor2_2
XANTENNA__16551__A3 _02479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16206_ _01796_ _01801_ _01804_ _02217_ _01679_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__o311a_1
X_13418_ net696 _07009_ _07291_ net504 vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__o211a_1
XANTENNA__12022__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17186_ _02490_ net77 _02727_ net1957 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[469\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_231_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14398_ game.CPU.applesa.ab.absxs.body_y\[70\] net953 vssd1 vssd1 vccd1 vccd1 _08272_
+ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_180_Right_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ _01749_ _01756_ _02143_ _02148_ _01645_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__o311a_1
XANTENNA__12573__B2 game.CPU.applesa.ab.absxs.body_y\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13349_ _06627_ _06641_ _06643_ _06642_ net508 net702 vssd1 vssd1 vccd1 vccd1 _07223_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16451__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19718__CLK clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15511__A1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16068_ _03234_ net269 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_295_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_255_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15019_ net1215 net1241 net820 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__and3_1
XANTENNA__15067__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17264__A1 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09065__A game.CPU.applesa.ab.absxs.body_y\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19827_ clknet_leaf_38_clk game.writer.tracker.next_frame\[422\] net1331 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[422\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_242_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12978__X _06852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10887__B2 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18378__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14078__B2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12203__B net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18742__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_320_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_316_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19868__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13825__A1 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19758_ clknet_leaf_26_clk game.writer.tracker.next_frame\[353\] net1312 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[353\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12628__A2 game.CPU.applesa.twoapples.absxs.next_head\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_223_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_242_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09511_ net1149 game.CPU.applesa.ab.absxs.body_y\[49\] vssd1 vssd1 vccd1 vccd1 _03754_
+ sky130_fd_sc_hd__or2_1
XANTENNA__10639__A1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18709_ clknet_leaf_50_clk _01126_ _00446_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[67\]
+ sky130_fd_sc_hd__dfrtp_4
X_19689_ clknet_leaf_34_clk game.writer.tracker.next_frame\[284\] net1320 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[284\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_223_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09442_ net1154 game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1 vssd1 vccd1
+ vccd1 _03685_ sky130_fd_sc_hd__xor2_1
XANTENNA__16775__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18892__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13589__B1 _07462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09373_ net1088 _03398_ net823 net900 _03615_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout244_A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16790__A3 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19559__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16527__B1 _02465_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13969__B game.CPU.applesa.ab.check_walls.above.walls\[83\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_352_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_306_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_331_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10272__C1 game.CPU.applesa.ab.YMAX\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09885__D _04127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12013__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14553__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11489__B _05331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13985__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17457__A _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1320_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16361__A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19398__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13108__A3 _06981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16080__B net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_A net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1206_X net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17255__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_342_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14069__A1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12888__X _06762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14069__B2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12113__B net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_180_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18288__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13277__C1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12619__A2 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17007__A1 _02497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09709_ net1084 game.CPU.applesa.ab.absxs.body_x\[23\] vssd1 vssd1 vccd1 vccd1 _03952_
+ sky130_fd_sc_hd__xor2_1
X_10981_ game.CPU.applesa.ab.absxs.body_x\[73\] net321 vssd1 vssd1 vccd1 vccd1 _04871_
+ sky130_fd_sc_hd__nand2_1
X_12720_ net872 net967 vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__nand2_2
XFILLER_0_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16766__B1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15143__C game.CPU.applesa.ab.check_walls.above.walls\[171\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_356_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_282_Right_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12651_ game.CPU.applesa.ab.absxs.body_x\[6\] net371 net367 game.CPU.applesa.ab.absxs.body_y\[7\]
+ _06453_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__a221o_1
XANTENNA__14241__A1 game.CPU.applesa.ab.absxs.body_y\[113\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16536__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16781__A3 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_178_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ net745 _05490_ _05489_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__a21bo_1
XANTENNA__14982__C game.CPU.applesa.ab.check_walls.above.walls\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19911__RESET_B net1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15370_ _08878_ _08897_ _08911_ _08909_ vssd1 vssd1 vccd1 vccd1 _08912_ sky130_fd_sc_hd__o31a_1
XANTENNA__11055__B2 game.CPU.applesa.ab.absxs.body_y\[106\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12582_ game.CPU.applesa.ab.absxs.body_x\[8\] net382 vssd1 vssd1 vccd1 vccd1 _06459_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__16255__B _08028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_324_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14321_ _03270_ net1048 _08190_ _08191_ _08194_ vssd1 vssd1 vccd1 vccd1 _08195_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_191_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11533_ net820 net260 net316 game.CPU.applesa.ab.check_walls.above.walls\[45\] vssd1
+ vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__a22o_1
XANTENNA__10802__B2 game.CPU.applesa.ab.absxs.body_y\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14056__A net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17040_ net67 _02678_ _02683_ net1729 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[367\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18615__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_312_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14252_ game.CPU.applesa.ab.absxs.body_y\[23\] net941 vssd1 vssd1 vccd1 vccd1 _08126_
+ sky130_fd_sc_hd__or2_1
X_11464_ game.CPU.applesa.ab.check_walls.above.walls\[17\] net771 vssd1 vssd1 vccd1
+ vccd1 _05353_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_311_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13203_ _07073_ _07074_ _07075_ _07076_ net496 net684 vssd1 vssd1 vccd1 vccd1 _07077_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10415_ _04338_ _04340_ game.CPU.randy.f1.state\[0\] vssd1 vssd1 vccd1 vccd1 _04561_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09420__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11395_ game.CPU.applesa.ab.check_walls.above.walls\[89\] net771 vssd1 vssd1 vccd1
+ vccd1 _05284_ sky130_fd_sc_hd__xor2_1
X_14183_ _03353_ net962 net941 _03352_ _08056_ vssd1 vssd1 vccd1 vccd1 _08057_ sky130_fd_sc_hd__a221o_1
XANTENNA__16271__A _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09420__B2 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13134_ game.writer.tracker.frame\[168\] game.writer.tracker.frame\[169\] net990
+ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10346_ _04505_ _04514_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__nor2_1
XFILLER_0_277_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18991_ net1197 _00217_ _00662_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18765__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13504__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ game.writer.tracker.frame\[212\] game.writer.tracker.frame\[213\] net1027
+ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_280_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ net655 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__inv_2
XANTENNA__10523__S _04632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10277_ _04374_ _04390_ _04459_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__o31a_1
XANTENNA__10318__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11522__A1_N net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17246__A1 _02275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ _05409_ _05410_ _05413_ _05414_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__or4_1
XFILLER_0_224_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17873_ net582 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__inv_2
XANTENNA__18198__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13834__S net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19612_ clknet_leaf_18_clk game.writer.tracker.next_frame\[207\] net1308 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[207\] sky130_fd_sc_hd__dfrtp_1
X_16824_ net173 _02520_ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__nor2_2
XANTENNA__15615__A game.CPU.applesa.ab.check_walls.above.walls\[82\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13807__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19543_ clknet_leaf_49_clk game.writer.tracker.next_frame\[138\] net1295 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[138\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_232_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16755_ _02404_ net64 _02587_ net1570 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[178\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_220_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19090__Q game.CPU.applesa.ab.check_walls.above.walls\[135\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13967_ net1070 _03475_ _03479_ net949 _07840_ vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__a221o_1
XFILLER_0_220_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15706_ game.CPU.applesa.ab.check_walls.above.walls\[152\] net269 vssd1 vssd1 vccd1
+ vccd1 _01718_ sky130_fd_sc_hd__nand2_1
X_19474_ clknet_leaf_19_clk game.writer.tracker.next_frame\[69\] net1335 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[69\] sky130_fd_sc_hd__dfrtp_1
X_12918_ net490 _06791_ _06790_ net227 vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_204_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16757__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_278_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16686_ _02460_ net62 _02562_ net1904 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[134\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15053__C game.CPU.applesa.ab.check_walls.above.walls\[81\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13898_ net1073 _03410_ game.CPU.applesa.ab.check_walls.above.walls\[57\] net884
+ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_347_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18425_ net610 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__inv_2
X_15637_ _03329_ net332 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__xnor2_1
X_12849_ _06721_ _06722_ net494 vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_291_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12974__A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19652__RESET_B net1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18356_ net596 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__inv_2
X_15568_ _01452_ _01584_ _01585_ _06545_ _03363_ vssd1 vssd1 vccd1 vccd1 game.writer.updater.update.next\[1\]
+ sky130_fd_sc_hd__o32a_1
X_17307_ net1847 net723 _02759_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[558\]
+ sky130_fd_sc_hd__and3_1
X_14519_ net1 _08392_ vssd1 vssd1 vccd1 vccd1 _08393_ sky130_fd_sc_hd__nand2_2
XFILLER_0_315_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18287_ net620 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
XANTENNA__10494__A _03197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15499_ _01449_ _01463_ _01490_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__o21bai_1
X_17238_ net154 _02428_ net79 _02740_ net1608 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[508\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19540__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_287_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11102__B net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17169_ _02465_ net73 _02723_ net1958 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[456\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_53_clk_X clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09991_ game.CPU.apple_location2\[0\] _04208_ _04209_ net1978 vssd1 vssd1 vccd1 vccd1
+ _01373_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_283_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload29_A clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19690__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ net1082 vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_244_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12214__A game.CPU.applesa.ab.check_walls.above.walls\[175\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_255_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_327_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_68_clk_X clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16996__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_193_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09523__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_223_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout361_A net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout459_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12482__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09425_ net1146 net798 vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__nand2_1
XANTENNA__19070__CLK net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_353_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_338_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout247_X net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_255_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16763__A3 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19393__RESET_B net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18638__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ net1155 _03486_ net780 net906 vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a22o_1
XFILLER_0_176_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16075__B net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09287_ net1083 game.CPU.applesa.ab.check_walls.above.walls\[83\] vssd1 vssd1 vccd1
+ vccd1 _03530_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1156_X net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16515__A3 _02456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10260__A2 _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout995_A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12108__B net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18788__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__A1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_344_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1323_X net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__B2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10200_ net1081 _04391_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__or2_1
XFILLER_0_293_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11947__B net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11180_ game.CPU.applesa.ab.absxs.body_y\[79\] net397 vssd1 vssd1 vccd1 vccd1 _05070_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__14323__B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ game.CPU.randy.f1.c1.count\[1\] _04325_ _04324_ _04323_ vssd1 vssd1 vccd1
+ vccd1 _04326_ sky130_fd_sc_hd__a211o_1
XFILLER_0_246_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17915__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_208_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15138__C net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17228__A1 _02413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09705__A2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _04233_ _04269_ _04235_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_351_Right_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14977__C game.CPU.applesa.ab.check_walls.above.walls\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14870_ _08655_ _08656_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[17\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10720__B1 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ net231 _07694_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__or2_1
XANTENNA__09469__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19413__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_230_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09469__B2 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_355_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16540_ net146 _02311_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13752_ _07624_ _07625_ net481 vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__mux2_1
X_10964_ _03285_ net545 vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__nand2_1
XANTENNA__13670__C1 net188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__B game.CPU.walls.rand_wall.input2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12703_ net966 _06571_ _06575_ _06567_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__a22o_1
X_16471_ net1709 _02420_ _02423_ net112 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[58\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12794__A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13683_ game.writer.tracker.frame\[449\] game.writer.tracker.frame\[451\] game.writer.tracker.frame\[452\]
+ game.writer.tracker.frame\[450\] net975 net1014 vssd1 vssd1 vccd1 vccd1 _07557_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_356_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10895_ _04792_ _04796_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__xnor2_1
X_18210_ net665 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__inv_2
X_15422_ _01449_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__inv_2
XANTENNA__15170__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19190_ clknet_leaf_46_clk net351 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.x_final\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_12634_ _06428_ _06459_ _06461_ _06462_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__or4_1
XANTENNA__19563__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13422__C1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_316_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18141_ net635 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__inv_2
XFILLER_0_344_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15353_ game.writer.updater.commands.count\[2\] _08889_ vssd1 vssd1 vccd1 vccd1 _08895_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__17164__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12565_ game.CPU.applesa.ab.absxs.body_x\[116\] net382 vssd1 vssd1 vccd1 vccd1 _06442_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_331_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14304_ game.CPU.applesa.ab.absxs.body_y\[28\] net868 net882 game.CPU.applesa.ab.absxs.body_x\[29\]
+ vssd1 vssd1 vccd1 vccd1 _08178_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11516_ net744 _05397_ _05401_ _05402_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a2111oi_1
X_18072_ net647 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__inv_2
XFILLER_0_297_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15284_ _08817_ _08829_ _08836_ _08815_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_123_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16911__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16272__Y _02278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ game.CPU.applesa.ab.absxs.body_x\[65\] net379 vssd1 vssd1 vccd1 vccd1 _06373_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_297_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12018__B net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17023_ _02362_ _02678_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__and2b_1
X_14235_ game.CPU.applesa.ab.absxs.body_y\[112\] net988 vssd1 vssd1 vccd1 vccd1 _08109_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_269_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11447_ game.CPU.applesa.ab.check_walls.above.walls\[73\] net771 vssd1 vssd1 vccd1
+ vccd1 _05336_ sky130_fd_sc_hd__xor2_1
XANTENNA__10539__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_20_Left_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_278_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_308_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09608__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11200__A1 game.CPU.applesa.ab.absxs.body_x\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14166_ _08028_ _08039_ vssd1 vssd1 vccd1 vccd1 _08040_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11378_ game.CPU.applesa.ab.check_walls.above.walls\[179\] net762 vssd1 vssd1 vccd1
+ vccd1 _05267_ sky130_fd_sc_hd__xor2_1
XANTENNA__11200__B2 game.CPU.applesa.ab.absxs.body_y\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14233__B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13117_ _06989_ _06990_ net482 vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__mux2_1
X_10329_ game.CPU.randy.f1.a1.count\[1\] game.CPU.randy.f1.a1.count\[0\] net740 vssd1
+ vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__and3_1
X_14097_ net945 net829 vssd1 vssd1 vccd1 vccd1 _07971_ sky130_fd_sc_hd__or2_1
X_18974_ net1201 _00198_ _00645_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12034__A game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17219__A1 _02391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13048_ _06860_ _06921_ net175 vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17925_ net613 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__inv_2
XFILLER_0_294_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_280_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12969__A net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1250 net1251 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11873__A game.CPU.applesa.ab.check_walls.above.walls\[140\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1261 game.CPU.bodymain1.Direction\[1\] vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__clkbuf_2
X_17856_ _03175_ _03177_ _03179_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__and3_1
XFILLER_0_294_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16978__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1272 net1273 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__clkbuf_2
Xfanout1283 net1293 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__clkbuf_4
Xfanout1294 net1297 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12688__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16807_ _02496_ net108 _02602_ net1578 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[215\]
+ sky130_fd_sc_hd__a22o_1
X_17787_ net758 game.CPU.applesa.normal1.counter_flip vssd1 vssd1 vccd1 vccd1 _01362_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_31_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14999_ net1223 net1255 game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1
+ vccd1 vccd1 _00216_ sky130_fd_sc_hd__and3_1
XFILLER_0_233_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14453__B2 game.CPU.applesa.ab.absxs.body_y\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_346_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19526_ clknet_leaf_22_clk game.writer.tracker.next_frame\[121\] net1342 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[121\] sky130_fd_sc_hd__dfrtp_1
X_16738_ net163 net68 net110 _02581_ net1540 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[167\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19906__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19457_ clknet_leaf_38_clk game.writer.tracker.next_frame\[52\] net1332 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[52\] sky130_fd_sc_hd__dfrtp_1
X_16669_ net2005 _02550_ _02552_ net127 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[127\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_313_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12908__S net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09210_ game.CPU.applesa.ab.check_walls.above.walls\[154\] vssd1 vssd1 vccd1 vccd1
+ _03459_ sky130_fd_sc_hd__inv_2
XANTENNA__15080__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18408_ net602 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19388_ clknet_leaf_9_clk _01394_ _00968_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.snake_head_x\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10936__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ game.CPU.applesa.ab.check_walls.above.walls\[24\] vssd1 vssd1 vccd1 vccd1
+ _03390_ sky130_fd_sc_hd__inv_2
X_18339_ net594 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__inv_2
XANTENNA__13964__B1 game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_350_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12209__A game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18391__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18930__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09632__A1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09632__B2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09072_ game.CPU.applesa.ab.absxs.body_y\[104\] vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__inv_2
XFILLER_0_288_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_250_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13739__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13811__S0 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout207_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09518__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09974_ net900 net1261 vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__nand2_1
XANTENNA__10950__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_256_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19436__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout743_A _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_48_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_357_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19574__RESET_B net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12455__B1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19586__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_196_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_357_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11007__B net536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15702__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout910_A net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout531_X net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1273_X net1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09408_ net1082 game.CPU.applesa.ab.check_walls.above.walls\[131\] vssd1 vssd1 vccd1
+ vccd1 _03651_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10680_ _04606_ _04615_ net754 vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_353_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_326_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_175_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09339_ net911 game.CPU.applesa.ab.absxs.body_x\[88\] _03327_ net1155 _03578_ vssd1
+ vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__a221o_1
XFILLER_0_152_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_350_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17146__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_303_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12119__A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_306_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12350_ _06226_ _06222_ _06221_ _06224_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__and4b_1
XFILLER_0_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ _05174_ _05182_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_214_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12281_ game.CPU.applesa.ab.check_walls.above.walls\[95\] net422 vssd1 vssd1 vccd1
+ vccd1 _06167_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11232_ game.CPU.applesa.ab.absxs.body_x\[14\] net409 vssd1 vssd1 vccd1 vccd1 _05122_
+ sky130_fd_sc_hd__xnor2_1
X_14020_ _07886_ _07887_ _07888_ _07893_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__a211o_1
XANTENNA__14380__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10581__B _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11163_ _03273_ net325 net535 _03342_ _05052_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__a221o_1
XANTENNA__11275__A2_N net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16121__A1 game.CPU.applesa.ab.check_walls.above.walls\[178\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ _03518_ game.CPU.applesa.twoapples.x_final\[3\] game.CPU.applesa.twoapples.start_enable
+ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_262_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16672__A2 _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_186_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11094_ game.CPU.applesa.ab.absxs.body_y\[59\] net399 vssd1 vssd1 vccd1 vccd1 _04984_
+ sky130_fd_sc_hd__xnor2_1
X_15971_ game.CPU.applesa.ab.absxs.body_x\[65\] net474 vssd1 vssd1 vccd1 vccd1 _01983_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__13384__S net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17710_ net1272 _04439_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_264_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15165__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14922_ _08658_ _08698_ vssd1 vssd1 vccd1 vccd1 _08699_ sky130_fd_sc_hd__or2_1
X_10045_ net1274 game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_128_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_303_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18690_ clknet_leaf_61_clk _01107_ _00427_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[32\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17216__A4 _02619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18803__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold60 game.CPU.applesa.ab.absxs.body_y\[1\] vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19929__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold71 net44 vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 game.writer.tracker.frame\[240\] vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ _08802_ net194 _03040_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__and3b_1
XFILLER_0_215_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14853_ net1626 _08645_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[10\]
+ sky130_fd_sc_hd__xor2_1
Xhold93 game.CPU.kyle.L1.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_349_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12301__B net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16975__A3 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13804_ game.writer.tracker.frame\[418\] net845 net838 game.writer.tracker.frame\[417\]
+ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__o22a_1
X_17572_ _04257_ net428 _02835_ _02995_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__a211o_1
X_14784_ net139 _08602_ _08603_ vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__and3_1
X_11996_ net825 net297 net291 game.CPU.applesa.ab.check_walls.above.walls\[30\] vssd1
+ vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__o22ai_1
XANTENNA__16267__Y _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19311_ net1163 _00035_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.out_random_2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_16523_ _02280_ net144 vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__nor2_2
XANTENNA__16708__B _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13735_ net508 _07604_ _07605_ _07608_ net227 vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_67_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15612__B net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_275_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10947_ game.CPU.applesa.ab.absxs.body_y\[30\] net541 vssd1 vssd1 vccd1 vccd1 _04837_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__18953__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16727__A3 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_217_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19242_ clknet_leaf_17_clk _00073_ _00880_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_16454_ net206 _02411_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__nor2_8
XFILLER_0_280_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13666_ net244 _07436_ _07438_ _07420_ net188 vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__o311a_1
XANTENNA__15935__B2 game.CPU.applesa.ab.check_walls.above.walls\[123\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10878_ game.CPU.applesa.ab.apple_possible\[6\] _04779_ vssd1 vssd1 vccd1 vccd1 _04780_
+ sky130_fd_sc_hd__and2_2
XANTENNA__12749__A1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14228__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15405_ _08935_ _01430_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__nor2_1
X_19173_ clknet_leaf_4_clk _01292_ _00835_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12617_ net1267 net384 _06229_ _06230_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__o211a_1
XFILLER_0_332_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17137__B1 _02713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16385_ game.writer.tracker.frame\[35\] net721 _02360_ vssd1 vssd1 vccd1 vccd1 _02361_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_139_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13597_ net278 _07470_ net246 vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__o21ai_2
XANTENNA__16283__X _02286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_314_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12844__S1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16724__A _02257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18124_ net577 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__inv_2
X_15336_ game.writer.updater.commands.mode\[2\] _03364_ game.writer.updater.commands.mode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08878_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_152_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12548_ game.CPU.applesa.ab.absxs.body_y\[22\] net518 vssd1 vssd1 vccd1 vccd1 _06425_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_170_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16443__B _02403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18055_ net653 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__inv_2
XANTENNA__18712__Q game.CPU.applesa.ab.absxs.body_x\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15267_ _08814_ _08822_ vssd1 vssd1 vccd1 vccd1 _08823_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12316__X _06202_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_2 _02179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ game.CPU.applesa.ab.absxs.body_x\[28\] net381 vssd1 vssd1 vccd1 vccd1 _06356_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__14244__A game.CPU.applesa.ab.absxs.body_x\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13174__A1 game.writer.tracker.frame\[449\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17006_ _02496_ net91 _02673_ net1589 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[343\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09378__B1 game.CPU.applesa.ab.check_walls.above.walls\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_300_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_269_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14218_ _08084_ _08087_ _08088_ _08091_ vssd1 vssd1 vccd1 vccd1 _08092_ sky130_fd_sc_hd__or4_2
XANTENNA__15059__B net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11587__B net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15198_ _00019_ _08764_ _08765_ _08767_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_78_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_286_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19459__CLK clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_228_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17555__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14149_ _07924_ _07926_ _07927_ _07821_ vssd1 vssd1 vccd1 vccd1 _08023_ sky130_fd_sc_hd__o31a_1
Xfanout509 net515 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09625__X _03868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_308_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18957_ net1200 _00210_ _00628_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12699__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19192__D net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15075__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17908_ net668 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__inv_2
X_09690_ net1092 game.CPU.applesa.ab.absxs.body_x\[6\] vssd1 vssd1 vccd1 vccd1 _03933_
+ sky130_fd_sc_hd__nand2_1
X_18888_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[18\] _00583_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[18\] sky130_fd_sc_hd__dfrtp_1
Xfanout1080 game.CPU.bad_collision vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__buf_8
Xfanout1091 game.CPU.applesa.ab.snake_head_x\[2\] vssd1 vssd1 vccd1 vccd1 net1091
+ sky130_fd_sc_hd__clkbuf_8
X_17839_ game.writer.updater.commands.count\[7\] _03165_ _03155_ vssd1 vssd1 vccd1
+ vccd1 _03167_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_240_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_324_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_233_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18386__A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_339_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_355_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19509_ clknet_leaf_14_clk game.writer.tracker.next_frame\[104\] net1282 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[104\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10947__A game.CPU.applesa.ab.absxs.body_y\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout157_A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_239_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11660__A1 _03385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_335_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_252_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16905__Y _02643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15654__A1_N game.CPU.applesa.ab.check_walls.above.walls\[164\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16193__X _02205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout324_A game.CPU.applesa.ab.absxs.next_head\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_335_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1066_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09124_ net1048 vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13977__B game.CPU.applesa.ab.check_walls.above.walls\[81\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17143__A3 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09055_ game.CPU.applesa.ab.absxs.body_y\[68\] vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11963__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_331_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout112_X net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14154__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_328_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold530 game.writer.tracker.frame\[256\] vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_303_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout693_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold541 game.CPU.randy.f1.a1.count\[8\] vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13260__S1 net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold552 game.CPU.walls.rand_wall.counter2\[1\] vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 game.writer.tracker.frame\[561\] vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13993__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold574 game.writer.tracker.frame\[18\] vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_275_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17300__B1 _02383_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold585 game.writer.tracker.frame\[156\] vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 game.writer.tracker.frame\[130\] vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1119_X net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_218_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09957_ net1146 _04186_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__and2_1
XANTENNA__19453__Q game.writer.tracker.frame\[48\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_A _03376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14601__B net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ _04103_ _04104_ _04108_ _03892_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__o31a_1
XFILLER_0_271_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12121__B net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18296__A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_339_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ net570 _05364_ _05737_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_352_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16528__B _02376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12979__A1 net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10801_ game.CPU.applesa.ab.absxs.body_y\[32\] _04696_ _04697_ game.CPU.applesa.ab.absxs.body_y\[28\]
+ vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__a22o_1
XANTENNA__09711__A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout913_X net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09844__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ net809 net301 _05665_ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_196_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14329__A game.CPU.applesa.ab.absxs.body_x\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09844__B2 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13520_ _07392_ _07393_ net285 vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10732_ game.CPU.applesa.ab.absxs.body_y\[23\] _04645_ _04652_ game.CPU.applesa.ab.absxs.body_y\[19\]
+ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__a22o_1
XANTENNA__15151__C game.CPU.applesa.ab.check_walls.above.walls\[179\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10576__B net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12573__A2_N net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13451_ net496 _07324_ _07323_ net230 vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__a211o_1
X_10663_ game.CPU.applesa.ab.absxs.body_x\[24\] _04695_ _04698_ game.CPU.applesa.ab.absxs.body_x\[20\]
+ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16544__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12402_ _03228_ game.CPU.applesa.twoapples.absxs.next_head\[3\] vssd1 vssd1 vccd1
+ vccd1 _06279_ sky130_fd_sc_hd__nor2_1
XFILLER_0_307_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16170_ game.CPU.applesa.ab.absxs.body_x\[34\] net466 net342 _03347_ _01624_ vssd1
+ vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a221o_1
XANTENNA__11403__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13382_ net247 _07194_ _07199_ net190 vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__a31o_1
XANTENNA__12600__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10594_ game.CPU.applesa.ab.absxs.body_x\[99\] net263 _04668_ net929 vssd1 vssd1
+ vccd1 vccd1 _01142_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_270_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15121_ net1207 net1233 game.CPU.applesa.ab.check_walls.above.walls\[149\] vssd1
+ vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__and3_1
XANTENNA__11954__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11688__A game.CPU.applesa.ab.check_walls.above.walls\[61\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12333_ net523 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.absxs.next_head\[5\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__19601__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12588__A2_N net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11040__X _04930_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13156__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_188_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__14353__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15052_ net1217 net1244 game.CPU.applesa.ab.check_walls.above.walls\[80\] vssd1 vssd1
+ vccd1 vccd1 _00274_ sky130_fd_sc_hd__and3_1
XANTENNA__09158__A game.CPU.applesa.ab.check_walls.above.walls\[50\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16893__A2 _02238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12264_ _06148_ _06149_ _06146_ _06147_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__a211o_1
XFILLER_0_266_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16550__Y _02480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14003_ net886 game.CPU.applesa.ab.check_walls.above.walls\[136\] _03455_ net947
+ vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11706__A2 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ _05097_ _05102_ _05103_ _05104_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__or4_2
X_19860_ clknet_leaf_20_clk game.writer.tracker.next_frame\[455\] net1317 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[455\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12195_ game.CPU.applesa.ab.check_walls.above.walls\[30\] net420 vssd1 vssd1 vccd1
+ vccd1 _06081_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_266_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_120_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19751__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18811_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[14\] _00548_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _03325_ net405 vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19791_ clknet_leaf_35_clk game.writer.tracker.next_frame\[386\] net1345 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[386\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15607__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14511__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_275_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10390__B2 net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15954_ game.CPU.applesa.ab.check_walls.above.walls\[30\] net442 vssd1 vssd1 vccd1
+ vccd1 _01966_ sky130_fd_sc_hd__xnor2_1
X_18742_ clknet_leaf_10_clk _01159_ _00479_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_11077_ game.CPU.applesa.ab.absxs.body_y\[41\] net542 vssd1 vssd1 vccd1 vccd1 _04967_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__13864__C1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_235_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12131__A2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _04234_ _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__nor2_1
X_14905_ net1153 _08424_ vssd1 vssd1 vccd1 vccd1 _08682_ sky130_fd_sc_hd__nand2_1
X_18673_ clknet_leaf_10_clk _01090_ _00410_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[103\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_188_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15885_ _03453_ net343 vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14408__A1 game.CPU.applesa.ab.absxs.body_x\[44\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_223_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15605__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14408__B2 game.CPU.applesa.ab.absxs.body_x\[47\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_199_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17070__A2 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17624_ game.CPU.kyle.L1.cnt_20ms\[13\] game.CPU.kyle.L1.cnt_20ms\[12\] _03027_ game.CPU.kyle.L1.cnt_20ms\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__a31o_1
XANTENNA__12419__B1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14836_ _08635_ _08636_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_230_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_337_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09621__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17555_ net1243 _02923_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__nand2_1
X_14767_ game.CPU.randy.counter1.count\[6\] game.CPU.randy.counter1.count\[4\] game.CPU.randy.counter1.count\[3\]
+ game.CPU.randy.counter1.count\[2\] vssd1 vssd1 vccd1 vccd1 _08588_ sky130_fd_sc_hd__or4_1
XANTENNA__09835__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ game.CPU.applesa.ab.check_walls.above.walls\[149\] net386 vssd1 vssd1 vccd1
+ vccd1 _05866_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_103_Left_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13631__A2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__B2 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16506_ net244 _02401_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__or2_1
XANTENNA__11215__X _05105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ game.writer.tracker.frame\[225\] game.writer.tracker.frame\[227\] game.writer.tracker.frame\[228\]
+ game.writer.tracker.frame\[226\] net968 net1000 vssd1 vssd1 vccd1 vccd1 _07592_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__19131__CLK net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17486_ _02910_ _02912_ _02914_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_329_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14698_ _08493_ _08495_ _08496_ _08536_ vssd1 vssd1 vccd1 vccd1 _08537_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16437_ game.writer.tracker.frame\[49\] _02395_ _02398_ net111 vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[49\] sky130_fd_sc_hd__a22o_1
X_19225_ clknet_leaf_66_clk _01319_ _00864_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_location\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13649_ net216 _07516_ net286 vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__o21a_1
XANTENNA__16454__A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16581__B2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13395__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09599__B1 game.CPU.applesa.ab.absxs.body_y\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_317_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14592__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19156_ clknet_leaf_70_clk _01277_ _00827_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.counter2\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_143_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16368_ net1997 net734 _02346_ _02349_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[29\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_309_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_288_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18107_ net632 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__inv_2
XANTENNA__19281__CLK clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15319_ game.CPU.applesa.twomode.number\[5\] _08859_ vssd1 vssd1 vccd1 vccd1 _08864_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19087_ net1178 _00124_ _00758_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[132\]
+ sky130_fd_sc_hd__dfrtp_1
X_16299_ net199 _02297_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__and2_4
XANTENNA__12046__X _05933_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18849__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18038_ net613 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__inv_2
XANTENNA__14344__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Left_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12206__B net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_319_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11110__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_300_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20000_ clknet_leaf_45_clk _01424_ net1300 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout306 net307 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16620__C _02375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09811_ net1155 game.CPU.applesa.ab.absxs.body_y\[24\] vssd1 vssd1 vccd1 vccd1 _04054_
+ sky130_fd_sc_hd__nand2_1
Xfanout317 net318 vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_4
Xfanout328 _04678_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_6
X_19989_ clknet_leaf_44_clk _01413_ net1305 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload11_A clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10381__B2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18999__CLK net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_302_Left_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09742_ net1140 net814 vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_253_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09673_ _03909_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__or2_1
XANTENNA__16188__X _02200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout274_A _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16939__A3 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13752__S net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11881__A1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_121_Left_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout441_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1183_A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10436__A2 _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_194_Right_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_311_Left_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1350_A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19624__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout706_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_323_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12808__S1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1069_X net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_323_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_350_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_323_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16083__B net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09107_ game.CPU.applesa.ab.absxs.body_y\[9\] vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__inv_2
XANTENNA__16514__D net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16324__A1 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_304_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1236_X net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_350_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16875__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19774__CLK clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_249_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_211_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09038_ game.CPU.applesa.ab.absxs.body_x\[117\] vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_300_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16370__Y _02351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11020__B net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold360 game.writer.tracker.frame\[510\] vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 game.writer.tracker.frame\[391\] vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 game.writer.tracker.frame\[277\] vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_276_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16088__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold393 game.writer.tracker.frame\[55\] vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _04883_ _04884_ _04885_ _04886_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a22o_1
XANTENNA__16627__A2 _02518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15427__B _01454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19004__CLK net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 _06598_ vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_183_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout851 _03494_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__buf_2
XFILLER_0_309_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09425__B net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout862 net863 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13846__C1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15146__C game.CPU.applesa.ab.check_walls.above.walls\[174\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout873 net875 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__buf_4
Xfanout884 net885 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_125_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13310__A1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09514__B1 game.CPU.applesa.ab.absxs.body_x\[48\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_300_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout895 net896 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_8
X_12951_ _06744_ _06746_ net676 vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__mux2_1
XANTENNA__10124__A1 net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_245_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11971__A game.CPU.applesa.ab.apple_possible\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__17052__A2 _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11902_ game.CPU.applesa.ab.check_walls.above.walls\[45\] net309 _05784_ _05788_
+ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__10675__A2 game.CPU.applesa.ab.absxs.body_x\[114\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15670_ game.CPU.applesa.ab.check_walls.above.walls\[107\] net458 vssd1 vssd1 vccd1
+ vccd1 _01682_ sky130_fd_sc_hd__nor2_1
XANTENNA__11872__A1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12882_ _06752_ _06753_ _06754_ _06755_ net481 net676 vssd1 vssd1 vccd1 vccd1 _06756_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_197_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14621_ game.CPU.clock1.counter\[12\] _08469_ net741 vssd1 vssd1 vccd1 vccd1 _08471_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__11690__B net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11833_ net789 net310 vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__or2_1
XANTENNA__10587__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09817__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_261_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09817__B2 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _08751_ _08753_ _02769_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12821__A0 _06690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14552_ net1175 game.CPU.walls.abc.number_out\[3\] vssd1 vssd1 vccd1 vccd1 _08421_
+ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_272_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11764_ net570 _05267_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13503_ net224 _07293_ _07376_ net274 vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__o211a_1
X_17271_ net112 _02489_ _02748_ net1921 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[533\]
+ sky130_fd_sc_hd__a22o_1
X_10715_ game.CPU.applesa.ab.absxs.body_y\[55\] _04609_ _04637_ game.CPU.applesa.ab.absxs.body_y\[51\]
+ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_342_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_194_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _08254_ _08258_ _08230_ vssd1 vssd1 vccd1 vccd1 _08357_ sky130_fd_sc_hd__a21oi_2
X_11695_ game.CPU.applesa.ab.check_walls.above.walls\[161\] net769 vssd1 vssd1 vccd1
+ vccd1 _05584_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19010_ net1189 _00238_ _00681_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[55\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_153_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16222_ net1447 _02232_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[0\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_82_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_341_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13434_ _06934_ _06937_ net702 vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_311_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ game.CPU.bad_collision _03244_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_12_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17107__A3 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16153_ _03459_ net347 net430 net788 _01717_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13365_ net479 _07238_ _07237_ net227 vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10577_ net936 net1266 _04657_ _04661_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__a31o_1
XFILLER_0_279_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15104_ net1204 net1231 net793 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ _06093_ _06094_ _06095_ _06166_ _06167_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__o32a_2
XANTENNA__16866__A2 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16084_ game.CPU.applesa.ab.check_walls.above.walls\[146\] net346 vssd1 vssd1 vccd1
+ vccd1 _02096_ sky130_fd_sc_hd__xnor2_1
X_13296_ _06775_ _06777_ net706 vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12026__B net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19912_ clknet_leaf_22_clk game.writer.tracker.next_frame\[507\] net1343 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[507\] sky130_fd_sc_hd__dfrtp_1
X_15035_ net1221 net1249 net816 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12247_ net798 net548 vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_283_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_286_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16618__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19843_ clknet_leaf_36_clk game.writer.tracker.next_frame\[438\] net1354 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[438\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_225_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09616__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11865__B net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ _06062_ _06063_ _06064_ _06058_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__o31a_1
XFILLER_0_219_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11129_ _03304_ net535 vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__xnor2_1
X_19774_ clknet_leaf_26_clk game.writer.tracker.next_frame\[369\] net1313 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[369\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_208_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_296_Right_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16986_ _02468_ net86 net715 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__o21a_1
X_18725_ clknet_leaf_63_clk _01142_ _00462_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[99\]
+ sky130_fd_sc_hd__dfrtp_4
X_15937_ _01940_ _01941_ _01942_ _01948_ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__or4_1
XANTENNA__16449__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13852__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17043__A2 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15868_ _01874_ _01875_ _01876_ _01878_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__or4_1
X_18656_ clknet_leaf_53_clk _01073_ _00393_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[70\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10666__A2 _04699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_305_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12696__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14819_ game.CPU.randy.counter1.count\[15\] _08624_ vssd1 vssd1 vccd1 vccd1 _08626_
+ sky130_fd_sc_hd__and2_1
X_17607_ _03020_ net429 _03019_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__and3b_1
XANTENNA__15072__B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19647__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18587_ clknet_leaf_31_clk _01007_ _00324_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[56\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_86_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09808__A1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10497__A _03197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15799_ game.CPU.applesa.ab.absxs.body_x\[50\] net467 net344 _03271_ vssd1 vssd1
+ vccd1 vccd1 _01811_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_294_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09808__B2 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_236_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17538_ net1273 _02829_ _02926_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__a21o_1
XANTENNA__09284__A2 _03527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_321_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17469_ _02889_ _02799_ _02894_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__mux2_1
XANTENNA__11105__B net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16554__A1 game.writer.tracker.frame\[81\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_190_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_345_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16554__B2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13601__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19208_ clknet_leaf_69_clk _00087_ _00856_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.YMAX\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18671__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19797__CLK clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_332_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10944__B net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload59_A clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__A2 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19139_ net1184 _00181_ _00810_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[184\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_298_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16857__A2 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_325_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_285_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18900__Q game.CPU.applesa.ab.good_collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13964__A1_N net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_247_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1029_A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16350__C _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout103 net110 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_285_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_273_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09526__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout114 _02243_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_8
XANTENNA__20004__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout125 net126 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout391_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 _02233_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout489_A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout147 net148 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_2
Xfanout158 net159 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_8
XANTENNA__17282__A2 _02258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19177__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout169 net170 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16490__B1 _02436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_263_Right_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09725_ net1081 _03231_ game.CPU.applesa.ab.absxs.body_x\[86\] net919 vssd1 vssd1
+ vccd1 vccd1 _03968_ sky130_fd_sc_hd__a22o_1
XANTENNA__16359__A net160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13843__A2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13335__X _07209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ net910 game.CPU.applesa.ab.check_walls.above.walls\[168\] game.CPU.applesa.ab.check_walls.above.walls\[169\]
+ net915 _03893_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__a221o_1
XANTENNA__10657__A2 _04696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_336_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09587_ _03826_ _03827_ _03828_ _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15550__X net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1186_X net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_328_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_258_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10200__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_231_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15710__B net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1353_X net1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16545__B2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10500_ net848 _04616_ _04622_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__or3_4
XFILLER_0_323_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11480_ game.CPU.applesa.ab.check_walls.above.walls\[48\] net777 vssd1 vssd1 vccd1
+ vccd1 _05369_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_323_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14326__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10431_ net1261 _04575_ _04573_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11302__Y game.CPU.applesa.ab.absxs.collision vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16381__X _02359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_208_Left_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_311_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12127__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14308__B1 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ game.writer.tracker.frame\[184\] game.writer.tracker.frame\[185\] net1039
+ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_304_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_347_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout980_X net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10362_ game.CPU.walls.rand_wall.input2 game.CPU.walls.rand_wall.counter2\[1\] game.CPU.walls.rand_wall.counter2\[0\]
+ game.CPU.walls.rand_wall.inputa vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__or4_1
XFILLER_0_289_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12319__C1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13657__S net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ net799 net555 vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11966__A _05731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13081_ _06947_ _06954_ net220 vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_269_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10293_ _03214_ net1442 _04473_ _04479_ vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout92_X net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15520__A2 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12414__X _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09436__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ game.CPU.applesa.ab.check_walls.above.walls\[141\] net386 vssd1 vssd1 vccd1
+ vccd1 _05919_ sky130_fd_sc_hd__xnor2_1
Xhold190 game.writer.tracker.frame\[504\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_256_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17273__A2 _02491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16840_ _02533_ net102 _02616_ net1607 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[234\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout670 _08799_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__buf_2
XANTENNA__14996__B net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout681 _06600_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_230_Right_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16771_ _02561_ _02592_ net736 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__o21a_1
XANTENNA__13295__A0 _06757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout692 _06600_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__buf_2
XFILLER_0_260_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_217_Left_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13983_ net1047 game.CPU.applesa.ab.check_walls.above.walls\[19\] vssd1 vssd1 vccd1
+ vccd1 _07857_ sky130_fd_sc_hd__or2_1
XANTENNA__16269__A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15722_ _03308_ net452 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__nand2_1
X_18510_ net579 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__inv_2
X_12934_ net211 _06708_ _06807_ net278 vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_358_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ clknet_leaf_23_clk game.writer.tracker.next_frame\[85\] net1339 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[85\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11845__B2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_220_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_358_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09171__A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18441_ net589 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__inv_2
X_15653_ net786 net430 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__xnor2_1
X_12865_ _06734_ _06735_ _06737_ _06736_ net476 net677 vssd1 vssd1 vccd1 vccd1 _06739_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_213_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14604_ game.CPU.clock1.counter\[5\] game.CPU.clock1.counter\[6\] _08458_ vssd1 vssd1
+ vccd1 vccd1 _08460_ sky130_fd_sc_hd__and3_1
XFILLER_0_157_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18372_ net598 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__inv_2
XANTENNA__18694__CLK clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11816_ net573 _05319_ _05320_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__a21oi_1
X_15584_ _01588_ _01589_ _01592_ _01593_ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__or4_1
X_12796_ game.writer.tracker.frame\[340\] game.writer.tracker.frame\[341\] net1029
+ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17323_ net1898 net732 _02763_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[570\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14535_ game.writer.control.current\[1\] _06547_ _08408_ game.writer.control.current\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08409_ sky130_fd_sc_hd__a31o_1
XFILLER_0_173_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11747_ _05632_ _05634_ _05626_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__and3b_1
XANTENNA__15620__B net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_299_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13421__A _06600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17254_ net175 _02287_ _02744_ net1806 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[520\]
+ sky130_fd_sc_hd__a22o_1
X_14466_ _03239_ net1066 net955 _03305_ _08339_ vssd1 vssd1 vccd1 vccd1 _08340_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_226_Left_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11678_ net816 net261 vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19088__Q game.CPU.applesa.ab.check_walls.above.walls\[133\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14236__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16205_ _02214_ _02215_ _02216_ _02213_ _02210_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__o311a_1
XANTENNA__16551__A4 _02480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13417_ net676 _07010_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__or2_1
XFILLER_0_342_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17185_ net149 _02327_ net77 _02727_ net1776 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[468\]
+ sky130_fd_sc_hd__a32o_1
X_10629_ _04682_ game.CPU.applesa.ab.absxs.body_x\[58\] net327 vssd1 vssd1 vccd1 vccd1
+ _01121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14397_ game.CPU.applesa.ab.absxs.body_y\[70\] net953 vssd1 vssd1 vccd1 vccd1 _08271_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_231_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13770__A1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16839__A2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16136_ _01768_ _02144_ _02145_ _02147_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__or4_4
X_13348_ _06620_ _06645_ _06646_ _06647_ net509 net703 vssd1 vssd1 vccd1 vccd1 _07222_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13567__S net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16067_ net780 net431 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__xnor2_1
X_13279_ game.writer.tracker.frame\[464\] game.writer.tracker.frame\[465\] net1013
+ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__mux2_1
XANTENNA__14252__A game.CPU.applesa.ab.absxs.body_y\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_295_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13522__A1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15018_ net1220 net1248 net821 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09346__A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11595__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_282_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11533__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19826_ clknet_leaf_38_clk game.writer.tracker.next_frame\[421\] net1329 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[421\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17264__A2 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_270_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_235_Left_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_320_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14078__A2 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09633__X _03876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_316_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19757_ clknet_leaf_26_clk game.writer.tracker.next_frame\[352\] net1312 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[352\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_223_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16969_ _02431_ net96 _02661_ net1826 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[318\]
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13825__A2 _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09510_ net1149 game.CPU.applesa.ab.absxs.body_y\[49\] vssd1 vssd1 vccd1 vccd1 _03753_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__15083__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17016__A2 net86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_242_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18708_ clknet_leaf_50_clk _01125_ _00445_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[66\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10639__A2 game.CPU.applesa.ab.absxs.body_x\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_19688_ clknet_leaf_34_clk game.writer.tracker.next_frame\[283\] net1320 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[283\] sky130_fd_sc_hd__dfrtp_1
X_09441_ _03678_ _03679_ _03681_ _03683_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__or4_2
XFILLER_0_91_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18639_ clknet_leaf_59_clk _01056_ _00376_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[37\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16775__A1 _02432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18394__A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_332_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_337_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10020__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09372_ net1130 game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1 vccd1
+ vccd1 _03615_ sky130_fd_sc_hd__xor2_1
XFILLER_0_176_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14250__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16527__B2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_305_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_331_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_321_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19599__RESET_B net1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16642__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout404_A net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1146_A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12564__A2 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_332_Right_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13985__B game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13477__S net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11786__A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1313_A net1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14162__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13513__A1 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_246_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18567__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19812__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17255__A2 _02466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_342_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1101_X net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_180_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout940_A game.CPU.applesa.y\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17007__A2 net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ net1130 game.CPU.applesa.ab.absxs.body_y\[23\] vssd1 vssd1 vccd1 vccd1 _03951_
+ sky130_fd_sc_hd__xor2_1
X_10980_ game.CPU.applesa.ab.absxs.body_x\[75\] net544 vssd1 vssd1 vccd1 vccd1 _04870_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_186_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19962__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09639_ net1145 _03461_ _03462_ net1135 _03881_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__a221o_1
XFILLER_0_356_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16766__A1 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_356_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12650_ _06274_ _06276_ _06480_ _06526_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__or4_1
XANTENNA__14241__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16536__B net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ game.CPU.applesa.ab.check_walls.above.walls\[98\] net768 vssd1 vssd1 vccd1
+ vccd1 _05490_ sky130_fd_sc_hd__xor2_2
XFILLER_0_356_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_178_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ game.CPU.applesa.ab.absxs.body_y\[23\] net364 vssd1 vssd1 vccd1 vccd1 _06458_
+ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14320_ _03340_ net993 net946 _03337_ vssd1 vssd1 vccd1 vccd1 _08194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_191_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11532_ net820 net260 net316 game.CPU.applesa.ab.check_walls.above.walls\[45\] vssd1
+ vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__o22ai_1
XANTENNA__10802__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17191__A1 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14056__B net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ game.CPU.applesa.ab.absxs.body_x\[22\] net878 net987 _03317_ _08118_ vssd1
+ vssd1 vccd1 vccd1 _08125_ sky130_fd_sc_hd__a221o_1
XFILLER_0_324_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19951__RESET_B net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ net744 _05350_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__nor2_1
XANTENNA__16552__A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13202_ game.writer.tracker.frame\[394\] game.writer.tracker.frame\[395\] net1020
+ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__mux2_1
XANTENNA__19342__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ _04360_ _04560_ _04554_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__o21a_1
X_14182_ game.CPU.applesa.ab.absxs.body_x\[18\] net1055 vssd1 vssd1 vccd1 vccd1 _08056_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__10566__A1 game.CPU.applesa.ab.absxs.body_x\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11394_ game.CPU.applesa.ab.check_walls.above.walls\[90\] net768 vssd1 vssd1 vccd1
+ vccd1 _05283_ sky130_fd_sc_hd__xor2_2
XANTENNA__16271__B _02275_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13387__S net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10566__B2 game.CPU.applesa.ab.absxs.body_x\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13133_ _07005_ _07006_ net482 vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__mux2_1
XANTENNA__15168__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11696__A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_267_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16151__C1 _02162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10345_ game.CPU.randy.f1.a1.count\[0\] net741 net1990 vssd1 vssd1 vccd1 vccd1 _04514_
+ sky130_fd_sc_hd__a21oi_1
X_18990_ net1197 _00216_ _00661_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[35\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13504__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09166__A game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13064_ game.writer.tracker.frame\[216\] game.writer.tracker.frame\[217\] net1015
+ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__mux2_1
X_17941_ net652 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_280_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10276_ net1169 _04463_ _04464_ _04468_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12304__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19492__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ _05899_ _05900_ _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__or3b_1
XANTENNA__17246__A2 _02448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17872_ net582 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__inv_2
X_19611_ clknet_leaf_18_clk game.writer.tracker.next_frame\[206\] net1310 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[206\] sky130_fd_sc_hd__dfrtp_1
X_16823_ game.writer.tracker.frame\[227\] _02606_ vssd1 vssd1 vccd1 vccd1 _02607_
+ sky130_fd_sc_hd__and2_1
XANTENNA__15615__B net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_232_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13807__A2 _07674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19542_ clknet_leaf_49_clk game.writer.tracker.next_frame\[137\] net1296 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[137\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11818__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16754_ _02398_ net63 _02587_ net1724 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[177\]
+ sky130_fd_sc_hd__a22o_1
X_13966_ net887 game.CPU.applesa.ab.check_walls.above.walls\[176\] _03477_ net1045
+ vssd1 vssd1 vccd1 vccd1 _07840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_232_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16206__B1 _02217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output33_A net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12917_ _06675_ _06676_ net683 vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__mux2_1
X_15705_ game.CPU.applesa.ab.check_walls.above.walls\[153\] net471 net465 game.CPU.applesa.ab.check_walls.above.walls\[154\]
+ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__o22a_1
X_19473_ clknet_leaf_19_clk game.writer.tracker.next_frame\[68\] net1335 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[68\] sky130_fd_sc_hd__dfrtp_1
X_16685_ _02267_ net62 _02562_ net1851 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[133\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_204_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16757__A1 _02405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13897_ net961 _03414_ _07768_ _07770_ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_278_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18424_ net626 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__inv_2
XFILLER_0_347_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12848_ game.writer.tracker.frame\[306\] game.writer.tracker.frame\[307\] net1028
+ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__mux2_1
X_15636_ _03330_ net336 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_83_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_291_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14518__Y _08392_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15567_ _03363_ _06545_ _08408_ _08412_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__and4_1
X_18355_ net594 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12779_ _06649_ _06650_ _06651_ _06652_ net493 net688 vssd1 vssd1 vccd1 vccd1 _06653_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_334_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_302_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14247__A game.CPU.applesa.ab.absxs.body_y\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17306_ net162 _02240_ _02394_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__or3_1
X_14518_ _08376_ _08381_ _08391_ vssd1 vssd1 vccd1 vccd1 _08392_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_124_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17182__A1 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15498_ _01470_ _01521_ _01512_ _01492_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__a2bb2o_2
X_18286_ net642 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_155_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17237_ net154 _02424_ net79 _02740_ net1637 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[507\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_303_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14449_ _08312_ _08313_ _08321_ _08322_ vssd1 vssd1 vccd1 vccd1 _08323_ sky130_fd_sc_hd__or4b_1
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16462__A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_302_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17168_ _02462_ net73 net558 vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19195__D net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16119_ game.CPU.applesa.ab.check_walls.above.walls\[177\] net475 net445 game.CPU.applesa.ab.check_walls.above.walls\[181\]
+ _02130_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a221o_1
XANTENNA__19835__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15078__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17099_ _02336_ net72 net736 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__o21a_1
X_09990_ game.CPU.apple_location2\[1\] _04208_ _04209_ net1448 vssd1 vssd1 vccd1 vccd1
+ _01374_ sky130_fd_sc_hd__a22o_1
XFILLER_0_268_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14299__A2 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15496__A1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15496__B2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ net1263 vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_243_Left_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_244_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12214__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18389__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_327_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17237__A2 _02424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17293__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19809_ clknet_leaf_40_clk game.writer.tracker.next_frame\[404\] net1357 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[404\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19985__CLK clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11014__A1_N game.CPU.applesa.ab.absxs.body_x\[54\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_208_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15799__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11809__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09523__B net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12230__A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19215__CLK net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16748__A1 _02394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16196__X _02208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_204_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout354_A net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09883__C1 _04125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1096_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ net924 game.CPU.applesa.ab.check_walls.above.walls\[115\] net797 net903 _03666_
+ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_252_Left_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16356__B _02340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_255_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_338_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18625__Q game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09355_ _03595_ _03596_ _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout142_X net142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14157__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1263_A game.CPU.applesa.clk_body vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout619_A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19365__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17173__A1 _02470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09286_ _03529_ _00291_ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_7_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13996__A net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10260__A3 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16920__A1 _02341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_X net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1149_X net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09402__A2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout890_A _03368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16091__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_344_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout988_A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_261_Left_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12405__A game.CPU.applesa.ab.absxs.body_x\[54\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1316_X net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13000__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_266_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10130_ game.CPU.randy.f1.c1.max_i\[1\] game.CPU.randy.f1.c1.count\[2\] vssd1 vssd1
+ vccd1 vccd1 _04325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_286_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18299__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_208_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17228__A2 _02720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10061_ _04216_ _04267_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__nor2_1
XANTENNA__13593__S0 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15716__A game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_234_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout943_X net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16987__A1 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_214_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10720__A1 game.CPU.applesa.ab.absxs.body_y\[46\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13820_ _07692_ _07693_ net499 vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_317_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15154__C game.CPU.applesa.ab.check_walls.above.walls\[182\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13751_ game.writer.tracker.frame\[137\] game.writer.tracker.frame\[139\] game.writer.tracker.frame\[140\]
+ game.writer.tracker.frame\[138\] net969 net991 vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_355_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16739__A1 _02370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__A2 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10963_ game.CPU.applesa.ab.absxs.body_x\[119\] net406 vssd1 vssd1 vccd1 vccd1 _04853_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16547__A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_253_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12702_ _06559_ _06572_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__or2_1
XANTENNA__14993__C game.CPU.applesa.ab.check_walls.above.walls\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16470_ net169 _02341_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__and2_4
X_13682_ game.writer.tracker.frame\[453\] game.writer.tracker.frame\[455\] game.writer.tracker.frame\[456\]
+ game.writer.tracker.frame\[454\] net975 net1015 vssd1 vssd1 vccd1 vccd1 _07556_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__19708__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10894_ _04793_ _04794_ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__and3_1
XANTENNA__14214__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15421_ game.writer.updater.commands.cmd_num\[1\] _01448_ _08934_ vssd1 vssd1 vccd1
+ vccd1 _01449_ sky130_fd_sc_hd__mux2_2
X_12633_ game.CPU.applesa.ab.absxs.body_x\[9\] net377 net519 game.CPU.applesa.ab.absxs.body_y\[10\]
+ _06460_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__a221o_1
XANTENNA__14067__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12139__X _06026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15352_ _08890_ _08893_ vssd1 vssd1 vccd1 vccd1 _08894_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18140_ net635 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__inv_2
X_12564_ game.CPU.applesa.ab.absxs.body_x\[118\] net372 net520 game.CPU.applesa.ab.absxs.body_y\[118\]
+ _06440_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__a221o_1
XANTENNA__17164__A1 _02456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16553__Y _02483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14303_ game.CPU.applesa.ab.absxs.body_y\[28\] net868 net861 game.CPU.applesa.ab.absxs.body_y\[29\]
+ _08174_ vssd1 vssd1 vccd1 vccd1 _08177_ sky130_fd_sc_hd__a221o_1
XFILLER_0_170_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11203__B net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11515_ net832 net253 _05398_ _04450_ _05403_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18071_ net647 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__inv_2
XANTENNA__19858__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18732__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15283_ _08824_ _08829_ _08812_ vssd1 vssd1 vccd1 vccd1 _08836_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_352_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16911__A1 _02322_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12495_ game.CPU.applesa.ab.absxs.body_y\[81\] net523 vssd1 vssd1 vccd1 vccd1 _06372_
+ sky130_fd_sc_hd__xnor2_1
X_17022_ net203 _02664_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__nor2_2
XANTENNA__13725__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14234_ game.CPU.applesa.ab.absxs.body_x\[115\] net1050 vssd1 vssd1 vccd1 vccd1 _08108_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__17097__B _02700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11446_ net745 _05332_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10539__A1 _03197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12933__C1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_312_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_308_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14165_ _08038_ _08029_ _08032_ vssd1 vssd1 vccd1 vccd1 _08039_ sky130_fd_sc_hd__or3b_1
XANTENNA__11200__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11377_ net743 _05265_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13116_ game.writer.tracker.frame\[138\] game.writer.tracker.frame\[139\] net991
+ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__mux2_1
XANTENNA__18882__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10328_ _04493_ _04504_ game.CPU.randy.f1.a1.count\[9\] net739 vssd1 vssd1 vccd1
+ vccd1 _01299_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_277_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14096_ net945 net829 vssd1 vssd1 vccd1 vccd1 _07970_ sky130_fd_sc_hd__nand2_1
X_18973_ net1198 _00187_ _00644_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_292_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13047_ net207 _06903_ _06920_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__o21ai_1
XANTENNA__17219__A2 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_237_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17924_ net591 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__inv_2
XFILLER_0_280_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10259_ net747 net742 _03370_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__a21o_1
XANTENNA__14530__A _08028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18002__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16427__B1 _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12161__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1240 net1241 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09624__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11873__B net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1251 net1255 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__buf_2
X_17855_ _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__inv_2
XFILLER_0_218_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1262 game.CPU.bodymain1.Direction\[1\] vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16978__A1 _02252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1273 game.CPU.luck1.Qa\[2\] vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__buf_2
Xfanout1284 net1286 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__clkbuf_4
X_16806_ _02492_ net108 _02602_ net1538 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[214\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13336__S0 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1295 net1296 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09486__A1_N net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12050__A net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17786_ game.CPU.applesa.good_collision2 _03492_ _03129_ game.CPU.applesa.twoapples.start_enable
+ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_31_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15064__C net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14453__A2 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14998_ net1223 net1251 game.CPU.applesa.ab.check_walls.above.walls\[26\] vssd1 vssd1
+ vccd1 vccd1 _00215_ sky130_fd_sc_hd__and3_1
XANTENNA__13110__C1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19525_ clknet_leaf_22_clk game.writer.tracker.next_frame\[120\] net1342 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[120\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16737_ _02369_ net61 _02581_ net1624 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[166\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_319_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13949_ net1043 game.CPU.applesa.ab.check_walls.above.walls\[131\] vssd1 vssd1 vccd1
+ vccd1 _07823_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_73_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__14385__A2_N net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_241_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_339_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19456_ clknet_leaf_39_clk game.writer.tracker.next_frame\[51\] net1332 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[51\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19388__CLK clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16668_ net168 net155 _02434_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__and3_1
XFILLER_0_313_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14205__A2 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15080__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18407_ net603 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__inv_2
XFILLER_0_201_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15619_ _03425_ net336 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19873__RESET_B net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13413__B1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19387_ clknet_leaf_3_clk _01393_ _00967_ vssd1 vssd1 vccd1 vccd1 game.CPU.bodymain1.main.score\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_16599_ net147 _02512_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ game.CPU.applesa.ab.check_walls.above.walls\[21\] vssd1 vssd1 vccd1 vccd1
+ _03389_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18338_ net594 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__inv_2
XANTENNA__17155__A1 _02435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13964__B2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09632__A2 game.CPU.applesa.ab.absxs.body_x\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_161_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_350_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16463__Y _02418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09071_ game.CPU.applesa.ab.absxs.body_y\[106\] vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11113__B net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12924__S net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16902__A1 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15705__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18269_ net647 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_288_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13716__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_287_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_250_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload41_A clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_330_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11727__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_330_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13811__S1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17458__A2 _02773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09518__B net1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_268_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09973_ net896 _04189_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_283_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13575__S0 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1011_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_283_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1109_A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09534__A game.CPU.applesa.ab.snake_head_x\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16969__A1 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout471_A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10702__A1 game.CPU.applesa.ab.absxs.body_y\[76\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10702__B2 game.CPU.applesa.ab.absxs.body_y\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13327__S0 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18605__CLK clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10399__B _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13101__C1 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_358_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09821__X _04064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout736_A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16367__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_196_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1099_X net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09407_ net1145 net792 vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18755__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout903_A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1266_X net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__A game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_175_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09338_ _03579_ _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__nand2_1
XANTENNA__17146__A1 _02419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_350_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10769__A1 game.CPU.applesa.ab.absxs.body_y\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_35_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12119__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_149_Left_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11023__B net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ game.CPU.randy.counter1.count1\[1\] vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_334_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_306_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13707__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11300_ _05148_ _05186_ _05189_ _05185_ _04907_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12280_ _06059_ _06060_ _06164_ _06165_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__or4_1
XANTENNA__09709__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_214_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout893_X net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11231_ _03319_ net405 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_293_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12135__A _03418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15149__C game.CPU.applesa.ab.check_walls.above.walls\[177\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_259_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11162_ _03341_ game.CPU.applesa.ab.absxs.next_head\[5\] vssd1 vssd1 vccd1 vccd1
+ _05052_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16121__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13665__S net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10113_ _04316_ game.CPU.applesa.apple_location2_n\[4\] _04311_ vssd1 vssd1 vccd1
+ vccd1 _01344_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13566__S0 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16672__A3 _02357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11093_ _03338_ net540 vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__nand2_1
X_15970_ _03335_ net337 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_186_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16409__B1 _02378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_158_Left_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09444__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10044_ _04247_ _04251_ _04242_ _04245_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__and4b_2
X_14921_ _08668_ _08696_ _08666_ vssd1 vssd1 vccd1 vccd1 _08698_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_303_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_264_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold50 _01311_ vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17082__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 net47 vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 game.CPU.applesa.ab.count_luck\[6\] vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
X_17640_ game.CPU.kyle.L1.cnt_500hz\[3\] _08801_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__or2_1
Xhold83 game.writer.tracker.frame\[110\] vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ _08645_ _08646_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.c1.innerCount\[9\]
+ sky130_fd_sc_hd__nor2_1
Xhold94 game.writer.tracker.frame\[486\] vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19530__CLK clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14435__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_348_Left_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13803_ game.writer.tracker.frame\[419\] net711 net674 game.writer.tracker.frame\[420\]
+ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__o22a_1
X_14783_ game.CPU.randy.counter1.count\[2\] game.CPU.randy.counter1.count\[1\] vssd1
+ vssd1 vccd1 vccd1 _08603_ sky130_fd_sc_hd__nand2_1
X_17571_ net426 _02841_ _02821_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__a21o_1
XANTENNA__13643__B1 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_187_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11995_ _05879_ _05880_ _05881_ _05878_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_55_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_348_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19310_ net1164 _00034_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.out_random_2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_16522_ net1738 _02457_ _02461_ net125 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[71\]
+ sky130_fd_sc_hd__a22o_1
X_13734_ net488 _07606_ _07607_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__and3_1
XANTENNA__16708__C _02328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_201_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10946_ game.CPU.applesa.ab.absxs.body_y\[28\] net533 vssd1 vssd1 vccd1 vccd1 _04836_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17385__A1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_275_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14509__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19241_ clknet_leaf_17_clk _00072_ _00879_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_344_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16453_ net242 _02265_ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__or2_2
X_13665_ _07531_ _07538_ net281 vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__mux2_1
XANTENNA__16564__X _02490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19680__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15935__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ game.CPU.applesa.ab.apple_possible\[4\] game.CPU.applesa.ab.apple_possible\[5\]
+ net760 vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_167_Left_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12749__A2 _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15404_ _01431_ _08939_ _08935_ game.writer.updater.commands.cmd_num\[4\] vssd1 vssd1
+ vccd1 vccd1 _01432_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13946__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ _06412_ _06492_ _06438_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__or3b_1
X_16384_ net1907 net720 _02360_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[34\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__13946__B2 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19172_ clknet_leaf_4_clk _01291_ _00834_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17137__A1 _02404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13596_ _07466_ _07469_ net227 vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_314_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11957__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15335_ game.writer.updater.commands.mode\[2\] _03364_ game.writer.updater.commands.mode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08877_ sky130_fd_sc_hd__nor3_2
X_18123_ net578 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12547_ _03249_ net371 vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_67_clk_X clknet_leaf_67_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14525__A _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_297_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_269_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_357_Left_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18054_ net653 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__inv_2
XANTENNA__09619__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15266_ _08813_ _01264_ vssd1 vssd1 vccd1 vccd1 _08822_ sky130_fd_sc_hd__nand2_1
X_12478_ game.CPU.applesa.ab.absxs.body_x\[29\] net375 net370 game.CPU.applesa.ab.absxs.body_x\[30\]
+ _06354_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__a221o_1
XANTENNA__19096__Q game.CPU.applesa.ab.check_walls.above.walls\[141\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_3 _02179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09378__A1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14244__B net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17005_ _02491_ net84 _02673_ net1603 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[342\]
+ sky130_fd_sc_hd__a22o_1
X_14217_ _08085_ _08086_ _08090_ _08083_ vssd1 vssd1 vccd1 vccd1 _08091_ sky130_fd_sc_hd__a211o_1
XFILLER_0_285_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09378__B2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11429_ game.CPU.applesa.ab.check_walls.above.walls\[29\] net317 vssd1 vssd1 vccd1
+ vccd1 _05318_ sky130_fd_sc_hd__or2_1
X_15197_ _00019_ _08766_ vssd1 vssd1 vccd1 vccd1 _08767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_286_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_238_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_300_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_238_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14148_ _07771_ _07776_ _07865_ _08021_ vssd1 vssd1 vccd1 vccd1 _08022_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_228_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14123__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_176_Left_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11884__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14123__B2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18956_ net1202 _00199_ _00627_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_14079_ net1172 net857 _07951_ _07952_ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__a22o_1
XANTENNA__18628__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12699__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17907_ net668 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__inv_2
XANTENNA__15075__B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18887_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[17\] _00582_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[17\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09550__A1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1070 net1071 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_206_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1081 net1083 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__buf_4
X_17838_ game.writer.updater.commands.count\[7\] _03165_ vssd1 vssd1 vccd1 vccd1 _03166_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09550__B2 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_175_Right_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1092 net1095 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_4
XFILLER_0_206_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16458__Y _02415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16820__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11108__B net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15803__B net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_221_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17769_ _03109_ _03120_ _03122_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_46_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
X_19508_ clknet_leaf_14_clk game.writer.tracker.next_frame\[103\] net1282 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[103\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15091__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_308_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_185_Left_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10947__B net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_239_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19439_ clknet_leaf_43_clk game.writer.tracker.next_frame\[34\] net1303 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[34\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11660__A2 _05194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_252_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_340_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11124__A game.CPU.applesa.ab.absxs.body_y\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09123_ net1057 vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout317_A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1059_A game.CPU.applesa.x\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09054_ game.CPU.applesa.ab.absxs.body_y\[70\] vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__inv_2
XANTENNA__10620__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_288_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14154__B _08027_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_328_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19403__CLK clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold520 game.writer.tracker.frame\[571\] vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_288_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_349_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout105_X net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold531 game.writer.tracker.frame\[74\] vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 game.writer.tracker.frame\[33\] vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1226_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12373__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_194_Left_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold553 game.writer.tracker.frame\[191\] vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11715__A3 _04441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold564 game.writer.tracker.frame\[285\] vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13993__B game.CPU.applesa.ab.check_walls.above.walls\[73\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold575 game.writer.tracker.frame\[190\] vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19734__Q game.writer.tracker.frame\[329\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold586 game.writer.tracker.frame\[23\] vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17300__B2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold597 game.writer.tracker.frame\[419\] vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13548__S0 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_263_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_256_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09956_ net1261 game.CPU.bodymain1.Direction\[0\] vssd1 vssd1 vccd1 vccd1 _04186_
+ sky130_fd_sc_hd__nand2b_1
XANTENNA__14170__A game.CPU.applesa.ab.absxs.body_y\[105\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__19553__CLK clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09887_ _03663_ _03664_ _03665_ _04129_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12402__B game.CPU.applesa.twoapples.absxs.next_head\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17064__B1 _02689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13625__A0 game.writer.tracker.frame\[305\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11018__B net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_339_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13073__X _06947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_352_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ game.CPU.applesa.ab.absxs.body_y\[33\] _04696_ _04697_ game.CPU.applesa.ab.absxs.body_y\[29\]
+ vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__a22o_1
X_11780_ net749 _05226_ net392 net810 _05666_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__a221o_1
XANTENNA__09711__B game.CPU.applesa.ab.absxs.body_y\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09844__A2 game.CPU.applesa.ab.absxs.body_x\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_338_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14329__B net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__Y _05194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10731_ game.CPU.applesa.ab.absxs.body_y\[28\] net330 _04714_ game.CPU.applesa.ab.absxs.body_y\[24\]
+ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout906_X net906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13450_ _07016_ _07033_ net704 vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17119__A1 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10662_ game.CPU.applesa.ab.absxs.body_x\[25\] _04695_ _04698_ game.CPU.applesa.ab.absxs.body_x\[21\]
+ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16544__B net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12401_ game.CPU.applesa.ab.absxs.body_x\[95\] net528 vssd1 vssd1 vccd1 vccd1 _06278_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11969__A game.CPU.applesa.ab.check_walls.above.walls\[148\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ net245 _07241_ _07251_ _07254_ net183 vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__a221o_1
XANTENNA__11403__A2 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10873__A game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10593_ _03228_ net263 vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__nor2_1
XFILLER_0_307_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11321__X _05210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15120_ net1207 net1230 net790 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__and3_1
XANTENNA__16878__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12332_ net1162 _04218_ _06211_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__a21o_1
XANTENNA__09439__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11688__B net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_188_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15051_ net1215 net1241 net811 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13787__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12263_ game.CPU.applesa.ab.check_walls.above.walls\[167\] net421 vssd1 vssd1 vccd1
+ vccd1 _06149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_259_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_277_Right_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12364__B1 game.CPU.applesa.twoapples.absxs.next_head\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14002_ net1062 game.CPU.applesa.ab.check_walls.above.walls\[137\] vssd1 vssd1 vccd1
+ vccd1 _07876_ sky130_fd_sc_hd__xor2_1
XANTENNA__14999__B net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11214_ _05093_ _05096_ _05098_ _05099_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__or4_1
X_12194_ _05878_ _06079_ _05880_ _05879_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__or4bb_1
Xoutput40 net40 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
X_18810_ clknet_leaf_73_clk game.CPU.clock1.next_counter\[13\] _00547_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.clock1.counter\[13\] sky130_fd_sc_hd__dfrtp_1
X_11145_ game.CPU.applesa.ab.absxs.body_y\[98\] net403 vssd1 vssd1 vccd1 vccd1 _05035_
+ sky130_fd_sc_hd__or2_1
X_19790_ clknet_leaf_35_clk game.writer.tracker.next_frame\[385\] net1345 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[385\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14080__A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12116__B1 _06002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13313__C1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09174__A game.CPU.applesa.ab.check_walls.above.walls\[80\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18741_ clknet_leaf_8_clk _01158_ _00478_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_15953_ game.CPU.applesa.ab.check_walls.above.walls\[27\] net462 vssd1 vssd1 vccd1
+ vccd1 _01965_ sky130_fd_sc_hd__and2_1
X_11076_ _03344_ net534 vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_262_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16559__X _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18920__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ net1090 _04232_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__nor2_1
X_14904_ net1153 _08424_ vssd1 vssd1 vccd1 vccd1 _08681_ sky130_fd_sc_hd__nor2_1
X_18672_ clknet_leaf_10_clk _01089_ _00409_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[102\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_203_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15884_ game.CPU.applesa.ab.check_walls.above.walls\[143\] net430 vssd1 vssd1 vccd1
+ vccd1 _01896_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_243_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14408__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09461__X _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17623_ net2038 _03028_ _03030_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_199_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15623__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14835_ game.CPU.randy.f1.c1.count\[3\] _08632_ _04332_ vssd1 vssd1 vccd1 vccd1 _08636_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_203_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14079__X _07953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12419__B2 game.CPU.applesa.ab.absxs.body_y\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_291_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_316_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09621__B game.CPU.applesa.ab.check_walls.above.walls\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17554_ _02819_ _02976_ _02977_ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__or4_1
X_14766_ game.CPU.randy.counter1.count\[7\] game.CPU.randy.counter1.count\[5\] game.CPU.randy.counter1.count\[1\]
+ net266 vssd1 vssd1 vccd1 vccd1 _08587_ sky130_fd_sc_hd__o31a_1
X_11978_ game.CPU.applesa.ab.check_walls.above.walls\[149\] net386 vssd1 vssd1 vccd1
+ vccd1 _05865_ sky130_fd_sc_hd__nand2_1
XFILLER_0_336_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14239__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16505_ net147 _02448_ _02449_ net189 vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a22o_4
X_13717_ game.writer.tracker.frame\[229\] game.writer.tracker.frame\[231\] game.writer.tracker.frame\[232\]
+ game.writer.tracker.frame\[230\] net968 net998 vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10929_ net537 vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__inv_2
XFILLER_0_329_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17485_ _02913_ _02905_ _02904_ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__mux2_1
X_14697_ _08529_ _08531_ _08534_ _08535_ vssd1 vssd1 vccd1 vccd1 _08536_ sky130_fd_sc_hd__o211a_1
XFILLER_0_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19224_ clknet_leaf_69_clk _01318_ _00863_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_location\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_16436_ net171 _02318_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__nor2_4
X_13648_ net495 _07519_ _07520_ _07521_ net230 vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__a311o_1
XANTENNA_clkbuf_leaf_32_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14041__B1 game.CPU.applesa.ab.check_walls.above.walls\[115\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14526__Y _08400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_317_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09599__A1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19426__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19155_ clknet_leaf_3_clk _00291_ _00826_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.inputa
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09599__B2 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16367_ net137 _02258_ _02348_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__and3_1
X_13579_ net222 _07448_ _07452_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_310_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_288_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10602__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18106_ net630 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__inv_2
X_15318_ _08863_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__inv_2
X_16298_ net206 net197 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__nand2_4
X_19086_ net1177 _00123_ _00757_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[131\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13778__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18037_ net606 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15249_ net587 _08808_ vssd1 vssd1 vccd1 vccd1 _08810_ sky130_fd_sc_hd__nor2_2
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16470__A net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_257_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_244_Right_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19576__CLK clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_285_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_319_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13158__X _07032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout307 _05606_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_4
X_09810_ _04047_ _04051_ _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__or3_1
XANTENNA__15086__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 _05213_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_2
XANTENNA__09771__B2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19988_ clknet_leaf_44_clk _01412_ net1304 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout329 _04672_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_238_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ net1095 game.CPU.applesa.ab.check_walls.above.walls\[66\] vssd1 vssd1 vccd1
+ vccd1 _03984_ sky130_fd_sc_hd__xor2_1
XANTENNA__09084__A game.CPU.applesa.ab.absxs.body_y\[72\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_253_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18939_ net1176 _00078_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number_out\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12222__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17046__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__A game.CPU.applesa.ab.absxs.body_x\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09672_ _03910_ _03911_ _03912_ _03914_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__a211o_1
XFILLER_0_253_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09812__A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_178_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11881__A2 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14280__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_194_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12830__A1 game.writer.tracker.frame\[289\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout434_A net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16364__B net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18633__Q game.CPU.applesa.ab.absxs.body_y\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_351_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1343_A net1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_220_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12594__B1 game.CPU.applesa.twoapples.absxs.next_head\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09106_ game.CPU.applesa.ab.absxs.body_y\[116\] vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__inv_2
XANTENNA__19919__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_304_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_211_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09037_ game.CPU.applesa.ab.absxs.body_x\[118\] vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16380__A net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1131_X net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_211_Right_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold350 game.writer.tracker.frame\[62\] vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 game.writer.tracker.frame\[316\] vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_229_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15708__B net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 game.writer.tracker.frame\[87\] vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_291_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold383 game.writer.tracker.frame\[564\] vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 game.writer.tracker.frame\[188\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout82_A _02690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout830 game.CPU.applesa.ab.check_walls.above.walls\[13\] vssd1 vssd1 vccd1 vccd1
+ net830 sky130_fd_sc_hd__clkbuf_4
Xfanout841 net842 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_4
XFILLER_0_244_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout852 net855 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_183_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09939_ net1118 net1120 vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__nand2_1
XANTENNA__16379__X _02357_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 net866 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__buf_4
XFILLER_0_309_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_245_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout874 net875 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__buf_4
Xfanout885 _03369_ vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09514__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12950_ net505 _06823_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__or2_1
XANTENNA__09514__B2 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout896 _03202_ vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__buf_4
XANTENNA__19905__RESET_B net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_300_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18100__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11901_ game.CPU.applesa.ab.check_walls.above.walls\[45\] net309 net394 game.CPU.applesa.ab.check_walls.above.walls\[44\]
+ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__17052__A3 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12881_ game.writer.tracker.frame\[42\] game.writer.tracker.frame\[43\] net992 vssd1
+ vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__mux2_1
XANTENNA__15599__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11872__A2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_325_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14620_ game.CPU.clock1.counter\[12\] _08469_ vssd1 vssd1 vccd1 vccd1 _08470_ sky130_fd_sc_hd__and2_1
X_11832_ net794 net299 _05712_ _05713_ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_197_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14271__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_318_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10587__B _04665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_261_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14551_ net468 vssd1 vssd1 vccd1 vccd1 game.CPU.walls.rand_wall.abduyd.next_wall\[2\]
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19449__CLK clknet_leaf_48_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11763_ _04442_ _05265_ _05650_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_272_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16555__A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_261_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_346_Right_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13502_ net482 _07290_ _07292_ net204 vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__a211o_1
X_10714_ game.CPU.applesa.ab.absxs.body_y\[60\] net425 _04713_ net934 vssd1 vssd1
+ vccd1 vccd1 _01067_ sky130_fd_sc_hd__a22o_1
X_17270_ _02275_ _02327_ _02748_ net1842 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[532\]
+ sky130_fd_sc_hd__a22o_1
X_14482_ _08351_ _08354_ _08129_ vssd1 vssd1 vccd1 vccd1 _08356_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_194_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ net786 net258 vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_342_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19288__D net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13433_ _06943_ _06957_ _06961_ _06960_ net501 net700 vssd1 vssd1 vccd1 vccd1 _07307_
+ sky130_fd_sc_hd__mux4_1
X_16221_ net556 net141 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__nor2_1
XANTENNA__14574__A1 net1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10645_ _04691_ game.CPU.applesa.ab.absxs.body_x\[43\] _04690_ vssd1 vssd1 vccd1
+ vccd1 _01114_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_311_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19599__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16152_ game.CPU.applesa.ab.check_walls.above.walls\[153\] net472 net430 net788 _01715_
+ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a221o_1
X_13364_ _06674_ _06676_ net701 vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__mux2_1
XANTENNA__09169__A game.CPU.applesa.ab.check_walls.above.walls\[68\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_341_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10576_ _03254_ net234 vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__nor2_1
XFILLER_0_341_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12307__B net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15103_ net1203 net1229 game.CPU.applesa.ab.check_walls.above.walls\[131\] vssd1
+ vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__and3_1
X_12315_ _06114_ _06115_ _06122_ _06128_ _06078_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__o2111a_1
X_16083_ _03458_ net342 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11211__B net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13295_ _06757_ _06776_ net704 vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_239_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16290__A _02274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19911_ clknet_leaf_22_clk game.writer.tracker.next_frame\[506\] net1343 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[506\] sky130_fd_sc_hd__dfrtp_1
X_15034_ net1222 net1250 game.CPU.applesa.ab.check_walls.above.walls\[62\] vssd1 vssd1
+ vccd1 vccd1 _00255_ sky130_fd_sc_hd__and3_1
X_12246_ game.CPU.applesa.ab.check_walls.above.walls\[182\] net419 vssd1 vssd1 vccd1
+ vccd1 _06132_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12888__A1 game.writer.tracker.frame\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_239_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15618__B net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_310_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_283_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17276__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17748__A_N _04255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19842_ clknet_leaf_36_clk game.writer.tracker.next_frame\[437\] net1353 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[437\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_294_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_286_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16618__A3 _02369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_225_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09616__B game.CPU.applesa.ab.check_walls.above.walls\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12177_ game.CPU.applesa.ab.check_walls.above.walls\[95\] net293 net288 net805 vssd1
+ vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_275_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11128_ _03284_ net415 vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__nand2_1
X_19773_ clknet_leaf_29_clk game.writer.tracker.next_frame\[368\] net1291 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[368\] sky130_fd_sc_hd__dfrtp_1
X_16985_ net149 _02466_ net89 _02666_ game.writer.tracker.frame\[329\] vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.next_frame\[329\] sky130_fd_sc_hd__a32o_1
XANTENNA__16289__X _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17291__A3 _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15193__X _00017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_322_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18724_ clknet_leaf_70_clk _01141_ _00461_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[98\]
+ sky130_fd_sc_hd__dfrtp_4
X_11059_ _04940_ _04941_ _04942_ _04944_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__or4_2
X_15936_ game.CPU.applesa.ab.check_walls.above.walls\[123\] net457 net465 game.CPU.applesa.ab.check_walls.above.walls\[122\]
+ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__18010__A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16449__B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_299_Left_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18655_ clknet_leaf_50_clk _01072_ _00392_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[69\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15867_ _01871_ _01872_ _01873_ _01877_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11863__A2 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20039__1363 vssd1 vssd1 vccd1 vccd1 _20039__1363/HI net1363 sky130_fd_sc_hd__conb_1
X_17606_ game.CPU.kyle.L1.cnt_20ms\[7\] game.CPU.kyle.L1.cnt_20ms\[6\] _03003_ vssd1
+ vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_235_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14818_ _08624_ _08625_ net138 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__and3b_1
XANTENNA__09351__B game.CPU.applesa.ab.absxs.body_x\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18586_ clknet_leaf_60_clk _01006_ _00323_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[51\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14262__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15798_ _03342_ net342 net446 game.CPU.applesa.ab.absxs.body_y\[49\] _01809_ vssd1
+ vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_86_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_294_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17537_ net846 _02852_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_28_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14749_ game.CPU.randy.counter1.count1\[15\] _08571_ vssd1 vssd1 vccd1 vccd1 _08574_
+ sky130_fd_sc_hd__or2_1
XANTENNA__16465__A net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_236_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_313_Right_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_317_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17468_ _02885_ _02894_ _02895_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__or3_1
XANTENNA__16554__A2 _02481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19549__Q game.writer.tracker.frame\[144\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19207_ clknet_leaf_70_clk _00086_ _00855_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.YMAX\[1\]
+ sky130_fd_sc_hd__dfstp_2
X_16419_ net198 _02385_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__and2_2
XANTENNA__13368__A2 _06690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_333_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17399_ _02826_ _02828_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12576__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19138_ net1188 _00180_ _00809_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[183\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17503__A1 game.CPU.luck1.Qa\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11121__B net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16857__A3 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19069_ net1185 _00104_ _00740_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[114\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_298_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_325_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10960__B net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_247_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13540__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout104 net105 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09526__B game.CPU.applesa.ab.check_walls.above.walls\[127\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout115 net118 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__buf_2
XFILLER_0_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12233__A net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout126 net129 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout137 _02233_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_169_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout148 _02270_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13828__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17282__A3 _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout159 _02269_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_4
XANTENNA_fanout384_A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15544__A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ net925 game.CPU.applesa.ab.absxs.body_x\[87\] game.CPU.applesa.ab.absxs.body_x\[85\]
+ net914 _03966_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__a221o_1
XANTENNA__16490__B2 _02273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18628__Q game.CPU.applesa.ab.absxs.body_y\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09655_ net1135 _03473_ _03474_ net1127 _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a221o_1
XANTENNA__17034__A3 _02634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout172_X net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16927__X _02650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout551_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16242__A1 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1293_A net1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_222_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_336_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout649_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_clk sky130_fd_sc_hd__clkbuf_8
X_09586_ net1086 game.CPU.applesa.ab.check_walls.above.walls\[19\] vssd1 vssd1 vccd1
+ vccd1 _03829_ sky130_fd_sc_hd__xor2_1
XFILLER_0_194_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16793__A2 net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16646__Y _02542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_328_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_258_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1081_X net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1179_X net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19741__CLK clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14005__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_231_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16094__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_324_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_351_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12567__B1 game.CPU.applesa.twoapples.absxs.next_head\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11312__A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13764__C1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ game.CPU.left_button.eD1.Q2 _04564_ _04569_ _04574_ vssd1 vssd1 vccd1 vccd1
+ _04575_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_351_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10042__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12127__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11031__B net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10042__B2 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14308__B2 game.CPU.applesa.ab.absxs.body_x\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10361_ net1937 game.CPU.walls.rand_wall.counter2\[0\] _04523_ vssd1 vssd1 vccd1
+ vccd1 _01278_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_347_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19891__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12319__B1 _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12100_ net798 net387 vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__or2_1
XANTENNA__11790__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_249_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11151__A2_N net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13080_ _06952_ _06953_ net478 vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__mux2_1
XANTENNA__09717__A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_269_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10292_ net851 game.CPU.applesa.ab.good_spot_next game.CPU.applesa.ab.apple_location\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__a21o_1
XFILLER_0_276_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout973_X net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15520__A3 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12031_ _05911_ _05917_ _05894_ _05902_ _05910_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__o2111a_1
XANTENNA__09735__A1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13531__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 game.writer.tracker.frame\[415\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09735__B2 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold191 game.writer.tracker.frame\[138\] vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout85_X net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10345__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13819__A0 game.writer.tracker.frame\[401\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_298_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_244_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout660 net661 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__buf_4
XFILLER_0_260_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout671 net672 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11982__A game.CPU.applesa.ab.check_walls.above.walls\[181\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14996__C game.CPU.applesa.ab.check_walls.above.walls\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout682 net692 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_4
X_16770_ net167 _02504_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__nand2_4
Xfanout693 net694 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_4
X_13982_ net1047 game.CPU.applesa.ab.check_walls.above.walls\[19\] vssd1 vssd1 vccd1
+ vccd1 _07856_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_109_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15721_ _03307_ net446 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__nand2_1
X_12933_ net494 _06806_ _06805_ net229 vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__o211a_1
XANTENNA__19271__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_358_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_220_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_358_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18440_ net588 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__inv_2
XANTENNA__13047__A1 net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15652_ net787 net438 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_319_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12864_ _06736_ _06737_ net500 vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16556__Y _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ net1892 _08458_ _08459_ vssd1 vssd1 vccd1 vccd1 game.CPU.clock1.next_counter\[5\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_185_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18371_ net596 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__inv_2
XANTENNA__11206__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11815_ net573 _05319_ _05321_ _04441_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__15901__B net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12795_ game.writer.tracker.frame\[344\] game.writer.tracker.frame\[345\] net1028
+ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15583_ game.CPU.applesa.ab.check_walls.above.walls\[91\] net460 net440 net805 _01590_
+ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__a221o_1
XFILLER_0_200_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17322_ net130 _02425_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14534_ net1080 net1 vssd1 vssd1 vccd1 vccd1 _08408_ sky130_fd_sc_hd__nand2_1
X_11746_ game.CPU.applesa.ab.check_walls.above.walls\[158\] net299 _05627_ _05631_
+ _05633_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_315_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_140_Left_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_315_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17253_ net204 net111 net68 _02744_ net1588 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[519\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16572__X _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14465_ game.CPU.applesa.ab.absxs.body_y\[60\] net993 vssd1 vssd1 vccd1 vccd1 _08339_
+ sky130_fd_sc_hd__xor2_1
X_11677_ _05549_ _05550_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__a21oi_2
XANTENNA__12558__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16204_ _01690_ _01691_ _01692_ _02122_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__or4b_1
X_13416_ _07011_ _07032_ net676 vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__mux2_1
X_10628_ net933 game.CPU.applesa.ab.absxs.body_x\[54\] vssd1 vssd1 vccd1 vccd1 _04682_
+ sky130_fd_sc_hd__and2_1
X_17184_ net157 _02322_ net71 net727 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__o31a_1
X_14396_ game.CPU.applesa.ab.absxs.body_y\[71\] net946 vssd1 vssd1 vccd1 vccd1 _08270_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12022__A2 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_231_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_330_Left_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13347_ _07217_ _07220_ net282 vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16135_ _01769_ _01770_ _01771_ _02146_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__or4_1
X_10559_ game.CPU.applesa.ab.absxs.body_x\[22\] _04645_ _04652_ game.CPU.applesa.ab.absxs.body_x\[18\]
+ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__a22o_1
XANTENNA__10584__A2 _04663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13507__C1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09627__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13278_ game.writer.tracker.frame\[460\] game.writer.tracker.frame\[461\] net1011
+ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__mux2_1
X_16066_ game.CPU.applesa.ab.check_walls.above.walls\[198\] _08429_ vssd1 vssd1 vccd1
+ vccd1 _02078_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_228_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12324__Y game.CPU.applesa.twoapples.absxs.next_head\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14252__B net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09726__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ net808 net422 vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__xnor2_1
X_15017_ net1220 net1249 game.CPU.applesa.ab.check_walls.above.walls\[45\] vssd1 vssd1
+ vccd1 vccd1 _00236_ sky130_fd_sc_hd__and3_1
XFILLER_0_295_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09346__B game.CPU.applesa.ab.absxs.body_y\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_267_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15067__C game.CPU.applesa.ab.check_walls.above.walls\[95\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15592__A1_N net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19825_ clknet_leaf_38_clk game.writer.tracker.next_frame\[420\] net1328 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[420\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_282_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09914__X _04156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17264__A3 _02479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19614__CLK clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13583__S net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19756_ clknet_leaf_25_clk game.writer.tracker.next_frame\[351\] net1319 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[351\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_251_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16968_ _02432_ _02636_ net729 vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__o21a_1
XANTENNA__14483__B1 _08230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18707_ clknet_leaf_50_clk _01124_ _00444_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[65\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09362__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_250_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_242_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15919_ _03448_ net350 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15083__B net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19687_ clknet_leaf_34_clk game.writer.tracker.next_frame\[282\] net1320 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[282\] sky130_fd_sc_hd__dfrtp_1
X_16899_ net200 net53 net92 _02641_ net1550 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[268\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__12500__B game.CPU.applesa.twoapples.absxs.next_head\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16224__A1 _08028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_182_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09440_ net1087 _03270_ game.CPU.applesa.ab.absxs.body_y\[58\] net905 _03682_ vssd1
+ vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__a221o_1
X_18638_ clknet_leaf_59_clk _01055_ _00375_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[36\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_149_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19764__CLK clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16775__A2 _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_332_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09371_ net1103 _03397_ _03400_ net1148 _03610_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__a221o_1
X_18569_ clknet_leaf_8_clk _00989_ _00306_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12927__S net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13171__X _07045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkload71_A clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12892__S0 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10955__B net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10272__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14427__B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_331_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout132_A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12013__A2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16642__B net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18911__Q game.CPU.applesa.enable_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09965__A1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10971__A net1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1041_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10575__A2 game.CPU.applesa.ab.absxs.body_x\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_320_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11786__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14162__B net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_246_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout599_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15826__X _01838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_301_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_357_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19568__RESET_B net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1306_A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_226_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19294__CLK clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_342_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout766_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13346__X _07220_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_180_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13277__A1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_241_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14474__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ net1160 _03413_ _03943_ _03949_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1296_X net1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_179_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11307__A game.CPU.applesa.ab.check_walls.above.walls\[71\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09638_ net925 game.CPU.applesa.ab.check_walls.above.walls\[155\] game.CPU.applesa.ab.check_walls.above.walls\[158\]
+ net902 vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_356_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16766__A2 _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_306_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_328_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11026__B net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16120__A2_N net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_242_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15721__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ net1100 _03236_ _03300_ net1139 _03811_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__a221o_2
XANTENNA__12837__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_356_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ game.CPU.applesa.ab.check_walls.above.walls\[99\] net763 vssd1 vssd1 vccd1
+ vccd1 _05489_ sky130_fd_sc_hd__xnor2_2
XANTENNA__16536__C _02386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ game.CPU.applesa.ab.absxs.body_x\[23\] net529 vssd1 vssd1 vccd1 vccd1 _06457_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_178_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_309_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11531_ _05411_ _05417_ _05418_ _05419_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__or4_1
XFILLER_0_147_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_191_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17191__A2 _02498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250_ _03249_ net1055 net963 _03316_ _08123_ vssd1 vssd1 vccd1 vccd1 _08124_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11462_ game.CPU.applesa.ab.check_walls.above.walls\[19\] net763 vssd1 vssd1 vccd1
+ vccd1 _05351_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19917__Q game.writer.tracker.frame\[512\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13201_ game.writer.tracker.frame\[398\] game.writer.tracker.frame\[399\] net1020
+ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__mux2_1
XANTENNA__16552__B _02318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ _04344_ _04559_ _04557_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ game.CPU.applesa.ab.absxs.body_x\[16\] net890 net864 game.CPU.applesa.ab.absxs.body_y\[17\]
+ _08054_ vssd1 vssd1 vccd1 vccd1 _08055_ sky130_fd_sc_hd__a221o_1
XFILLER_0_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10881__A game.CPU.applesa.ab.apple_possible\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11393_ game.CPU.applesa.ab.check_walls.above.walls\[91\] net763 vssd1 vssd1 vccd1
+ vccd1 _05282_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10566__A2 _04653_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11763__A1 _04442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ _07002_ _07004_ net679 vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__mux2_1
X_20038__1362 vssd1 vssd1 vccd1 vccd1 _20038__1362/HI net1362 sky130_fd_sc_hd__conb_1
X_10344_ net740 _04488_ _04513_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_277_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_267_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19637__CLK clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13063_ game.writer.tracker.frame\[246\] game.writer.tracker.frame\[247\] net1030
+ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17940_ net640 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__inv_2
XFILLER_0_277_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_267_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10275_ net1172 _04375_ _04466_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_115_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_280_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19920__RESET_B net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11515__A1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ net811 net298 net290 net812 vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__o22a_1
XANTENNA__11515__B2 _04450_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17871_ _03367_ _03189_ _03184_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_292_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10105__B game.CPU.applesa.enable_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19610_ clknet_leaf_18_clk game.writer.tracker.next_frame\[205\] net1310 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[205\] sky130_fd_sc_hd__dfrtp_1
X_16822_ net131 net66 net122 _02606_ net1508 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[226\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__13268__A1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout490 net494 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_4
XANTENNA__18661__CLK clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19787__CLK clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19541_ clknet_leaf_33_clk game.writer.tracker.next_frame\[136\] net1301 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[136\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_232_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16753_ _02535_ _02561_ net735 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__o21a_1
X_13965_ net882 game.CPU.applesa.ab.check_walls.above.walls\[177\] game.CPU.applesa.ab.check_walls.above.walls\[181\]
+ net862 _07838_ vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__a221o_1
XANTENNA__18495__A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_260_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_232_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15704_ _03460_ net343 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__xnor2_1
X_19472_ clknet_leaf_19_clk game.writer.tracker.next_frame\[67\] net1335 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[67\] sky130_fd_sc_hd__dfrtp_1
X_12916_ net503 _06789_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__or2_1
XFILLER_0_220_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16684_ _02454_ net62 _02562_ net1894 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[132\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16757__A2 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_216_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_204_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09892__B1 _03737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ net870 net817 game.CPU.applesa.ab.check_walls.above.walls\[62\] net854 _07769_
+ vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__a221o_1
X_18423_ net626 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__inv_2
XANTENNA_output26_A net1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15635_ game.CPU.applesa.ab.absxs.body_x\[83\] net457 vssd1 vssd1 vccd1 vccd1 _01647_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12847_ game.writer.tracker.frame\[310\] game.writer.tracker.frame\[311\] net1033
+ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__mux2_1
XANTENNA__12779__A0 _06649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_347_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_291_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ net595 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__inv_2
X_15566_ _03363_ _01580_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_25_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ game.writer.tracker.frame\[122\] game.writer.tracker.frame\[123\] net1033
+ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__mux2_1
XANTENNA__16509__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14247__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17305_ net175 net116 _02390_ _02758_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[557\]
+ sky130_fd_sc_hd__a31o_1
X_14517_ _08388_ _08389_ _08390_ vssd1 vssd1 vccd1 vccd1 _08391_ sky130_fd_sc_hd__or3_2
XFILLER_0_327_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11729_ _05601_ _05602_ _05616_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__and3_1
X_18285_ net641 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
X_15497_ _06557_ _01508_ _01518_ _01520_ _01469_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_299_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17182__A2 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_315_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17236_ net157 _02425_ net72 net729 vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__o31a_1
XFILLER_0_114_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14448_ game.CPU.applesa.ab.absxs.body_y\[89\] net861 net949 _03326_ vssd1 vssd1
+ vccd1 vccd1 _08322_ sky130_fd_sc_hd__o22a_1
XFILLER_0_141_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11887__A game.CPU.applesa.ab.check_walls.above.walls\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_17167_ _02461_ net77 _02722_ net1774 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[455\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10892__D_N net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14379_ game.CPU.applesa.ab.absxs.body_y\[80\] net983 vssd1 vssd1 vccd1 vccd1 _08253_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11754__A1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_268_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11754__B2 game.CPU.applesa.ab.check_walls.above.walls\[173\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16118_ net783 net437 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15078__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16142__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17098_ net160 net69 net80 _02701_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[407\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_255_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16693__A1 _02300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08940_ net1080 vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__inv_2
X_16049_ game.CPU.applesa.ab.absxs.body_y\[103\] net432 vssd1 vssd1 vccd1 vccd1 _02061_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_244_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17293__B _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17237__A3 net79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_327_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15806__B net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_208_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_166_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19808_ clknet_leaf_37_clk game.writer.tracker.next_frame\[403\] net1354 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[403\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16996__A2 net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19739_ clknet_leaf_18_clk game.writer.tracker.next_frame\[334\] net1289 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[334\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11809__A2 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12230__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_343_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11127__A game.CPU.applesa.ab.absxs.body_x\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10031__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16748__A2 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12482__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14208__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09423_ net1107 game.CPU.applesa.ab.check_walls.above.walls\[112\] vssd1 vssd1 vccd1
+ vccd1 _03666_ sky130_fd_sc_hd__xor2_1
XFILLER_0_176_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10966__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_A game.CPU.walls.rand_wall.abduyd.next_wall\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_353_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_255_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09354_ net1085 _03289_ _03356_ net1149 vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1089_A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12865__S0 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10685__B net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14157__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17749__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ game.CPU.walls.rand_wall.count1 net756 _03527_ net755 vssd1 vssd1 vccd1 vccd1
+ _00291_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout514_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout135_X net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10796__A2 _04690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1256_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13996__B net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16920__A2 _02643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16372__B net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_278_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14173__A game.CPU.applesa.ab.absxs.body_y\[106\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_X net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11745__A1 game.CPU.applesa.ab.check_walls.above.walls\[156\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_344_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16133__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout883_A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16684__A1 _02454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_189_Right_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_266_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1211_X net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14901__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18684__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_208_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ _04236_ _04267_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_237_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15716__B net441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_274_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14447__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16987__A2 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10720__A2 _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_254_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_317_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_253_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15732__A game.CPU.applesa.ab.absxs.body_y\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_97_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13750_ game.writer.tracker.frame\[141\] game.writer.tracker.frame\[143\] game.writer.tracker.frame\[144\]
+ game.writer.tracker.frame\[142\] net966 net990 vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__mux4_1
X_10962_ game.CPU.applesa.ab.absxs.body_y\[119\] net398 vssd1 vssd1 vccd1 vccd1 _04852_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_355_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16739__A2 _02561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13670__B2 _07471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16547__B net146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ _06572_ net841 vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__nand2_1
XFILLER_0_329_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13681_ net221 _07548_ net284 vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__o21a_1
X_10893_ game.CPU.applesa.ab.XMAX\[0\] net773 _04449_ _04454_ vssd1 vssd1 vccd1 vccd1
+ _04795_ sky130_fd_sc_hd__a211o_1
XANTENNA__10876__A game.CPU.applesa.ab.apple_possible\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_195_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14348__A game.CPU.applesa.ab.absxs.body_x\[34\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_210_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11324__X _05213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15420_ _01445_ _01447_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_356_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_219_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12632_ _03290_ game.CPU.applesa.twoapples.absxs.next_head\[2\] net524 game.CPU.applesa.ab.absxs.body_y\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__a22o_1
XANTENNA__13422__A1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_195_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14067__B game.CPU.applesa.ab.check_walls.above.walls\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15351_ game.writer.updater.commands.count\[16\] game.writer.updater.commands.count\[12\]
+ _08891_ _08892_ vssd1 vssd1 vccd1 vccd1 _08893_ sky130_fd_sc_hd__or4_1
X_12563_ game.CPU.applesa.ab.absxs.body_x\[119\] net530 vssd1 vssd1 vccd1 vccd1 _06440_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_309_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17164__A2 _02720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16563__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_202_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14302_ game.CPU.applesa.ab.absxs.body_y\[31\] net939 vssd1 vssd1 vccd1 vccd1 _08176_
+ sky130_fd_sc_hd__xor2_1
X_11514_ net567 _05399_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18070_ net647 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__inv_2
X_12494_ game.CPU.applesa.ab.absxs.body_x\[81\] net375 net364 game.CPU.applesa.ab.absxs.body_y\[83\]
+ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__a2bb2o_1
X_15282_ _08815_ _08830_ _08835_ _08812_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_324_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16911__A2 _02636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19296__D net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13398__S net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17021_ net66 net85 _02677_ net1509 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[354\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09929__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14233_ game.CPU.applesa.ab.absxs.body_x\[112\] net1074 vssd1 vssd1 vccd1 vccd1 _08107_
+ sky130_fd_sc_hd__xor2_1
X_11445_ net745 _05332_ _05333_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14083__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10539__A2 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ net1131 net859 _08033_ _08035_ _08037_ vssd1 vssd1 vccd1 vccd1 _08038_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16124__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11376_ game.CPU.applesa.ab.check_walls.above.walls\[178\] net767 vssd1 vssd1 vccd1
+ vccd1 _05265_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_308_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13115_ game.writer.tracker.frame\[142\] game.writer.tracker.frame\[143\] net990
+ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ game.CPU.randy.f1.a1.count\[9\] _04491_ _04487_ vssd1 vssd1 vccd1 vccd1 _04504_
+ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14095_ net1068 _03383_ _03384_ net986 _07968_ vssd1 vssd1 vccd1 vccd1 _07969_ sky130_fd_sc_hd__a221o_1
X_18972_ net1199 _00176_ _00643_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13046_ net245 _06907_ _06911_ _06919_ net225 vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__a311o_1
X_17923_ net605 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__inv_2
XANTENNA__17219__A3 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10258_ net774 net769 vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__or2_2
XANTENNA__15626__B net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12161__A1 game.CPU.applesa.ab.check_walls.above.walls\[39\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16427__A1 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1230 net1231 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_2
Xfanout1241 net1242 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12161__B2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17854_ game.writer.updater.commands.count\[11\] game.writer.updater.commands.count\[10\]
+ _03169_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__and3_1
XFILLER_0_218_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09624__B game.CPU.applesa.ab.check_walls.above.walls\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_294_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1252 net1254 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__clkbuf_2
X_10189_ net1105 _04381_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__or2_1
XANTENNA__12331__A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16978__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1263 game.CPU.applesa.clk_body vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__buf_4
Xfanout1274 game.CPU.kyle.L1.row_2\[72\] vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__clkbuf_4
X_16805_ _02490_ net108 _02602_ net1739 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[213\]
+ sky130_fd_sc_hd__a22o_1
Xfanout1285 net1286 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13336__S1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1296 net1297 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__clkbuf_4
X_17785_ _03358_ _03128_ _03132_ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_227_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12050__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14997_ net1223 net1251 game.CPU.applesa.ab.check_walls.above.walls\[25\] vssd1 vssd1
+ vccd1 vccd1 _00214_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_31_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19524_ clknet_leaf_21_clk game.writer.tracker.next_frame\[119\] net1336 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[119\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15642__A game.CPU.applesa.ab.check_walls.above.walls\[73\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16736_ net184 _02524_ net101 _02581_ net1585 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[165\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_163_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13948_ net938 game.CPU.applesa.ab.check_walls.above.walls\[135\] vssd1 vssd1 vccd1
+ vccd1 _07822_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_319_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09640__A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19455_ clknet_leaf_39_clk game.writer.tracker.next_frame\[50\] net1332 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[50\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16667_ net1901 _02550_ _02551_ net127 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[126\]
+ sky130_fd_sc_hd__a22o_1
X_13879_ net877 game.CPU.applesa.ab.check_walls.above.walls\[106\] game.CPU.applesa.ab.check_walls.above.walls\[104\]
+ net887 vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14258__A game.CPU.applesa.ab.absxs.body_y\[79\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_234_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18406_ net603 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
XFILLER_0_243_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15618_ _03424_ net353 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13413__A1 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19386_ clknet_leaf_3_clk _01392_ _00966_ vssd1 vssd1 vccd1 vccd1 game.CPU.bodymain1.main.score\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_16598_ net167 _02437_ _02358_ _01516_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__18557__CLK clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18337_ net593 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15549_ _01540_ _01562_ _01569_ _01470_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_84_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19802__CLK clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09070_ game.CPU.applesa.ab.absxs.body_y\[13\] vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__inv_2
X_18268_ net648 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
XANTENNA__16902__A2 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17219_ _02391_ net122 net119 _02735_ net1495 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[494\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15089__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_250_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14913__A1 game.CPU.applesa.ab.XMAX\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19842__RESET_B net1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14913__B2 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18199_ net580 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
XANTENNA__11727__B2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_303_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_287_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19952__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload34_A clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_338_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12940__S net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09972_ net1136 net850 _04200_ vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_268_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_256_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10950__A2 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_228_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14440__B net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout297_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12241__A game.CPU.applesa.ab.check_walls.above.walls\[151\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09534__B game.CPU.applesa.ab.check_walls.above.walls\[74\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1004_A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16969__A2 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_271_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10702__A2 _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17091__A1 _02484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13327__S1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_224_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19332__CLK clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12455__A2 game.CPU.applesa.twoapples.absxs.next_head\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16367__B _02258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18636__Q game.CPU.applesa.ab.absxs.body_y\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10466__A1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_211_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout252_X net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09406_ net1089 game.CPU.applesa.ab.check_walls.above.walls\[130\] vssd1 vssd1 vccd1
+ vccd1 _03649_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_45_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_303_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19482__CLK clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09337_ net1098 game.CPU.applesa.ab.absxs.body_x\[89\] vssd1 vssd1 vccd1 vccd1 _03580_
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_258_Right_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_175_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1161_X net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_350_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10769__A2 _04675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ game.CPU.randy.counter1.count\[1\] vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09199_ game.CPU.applesa.ab.check_walls.above.walls\[129\] vssd1 vssd1 vccd1 vccd1
+ _03448_ sky130_fd_sc_hd__inv_2
XANTENNA__09709__B game.CPU.applesa.ab.absxs.body_x\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13011__S net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_214_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ game.CPU.applesa.ab.absxs.body_y\[15\] net398 vssd1 vssd1 vccd1 vccd1 _05120_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__11320__A game.CPU.applesa.ab.apple_possible\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_160_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_321_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_278_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14380__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16830__B _02524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12135__B net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16657__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_248_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11161_ _05045_ _05046_ _05048_ _05049_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a22o_1
XFILLER_0_219_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10112_ game.CPU.applesa.enable_in game.CPU.applesa.twoapples.y_final\[0\] _03212_
+ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__a21o_1
XFILLER_0_274_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13566__S1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_207_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11092_ game.CPU.applesa.ab.absxs.body_y\[58\] net401 vssd1 vssd1 vccd1 vccd1 _04982_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_186_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_274_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13340__B1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16409__B2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_234_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10043_ net1174 _04226_ _04249_ _04250_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__a22o_1
X_14920_ _08668_ _08696_ vssd1 vssd1 vccd1 vccd1 _08697_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09444__B game.CPU.applesa.ab.check_walls.above.walls\[143\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12151__A net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_303_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold40 game.CPU.applesa.twomode.number\[1\] vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17082__A1 _02303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold51 game.CPU.applesa.ab.y_final\[2\] vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 game.writer.tracker.frame\[0\] vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 game.CPU.applesa.ab.apple_location\[7\] vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ net1983 _08643_ vssd1 vssd1 vccd1 vccd1 _08646_ sky130_fd_sc_hd__nor2_1
Xhold84 game.writer.tracker.frame\[416\] vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_270_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold95 game.writer.tracker.frame\[239\] vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13802_ game.writer.tracker.frame\[422\] net845 net838 game.writer.tracker.frame\[421\]
+ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__o22a_1
X_17570_ net739 _02851_ _02950_ _02849_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__a22o_1
X_14782_ game.CPU.randy.counter1.count\[2\] game.CPU.randy.counter1.count\[1\] vssd1
+ vssd1 vccd1 vccd1 _08602_ sky130_fd_sc_hd__or2_1
X_11994_ game.CPU.applesa.ab.check_walls.above.walls\[29\] net388 vssd1 vssd1 vccd1
+ vccd1 _05881_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13643__B2 game.writer.tracker.frame\[32\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16521_ net212 net154 _02373_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__and3_2
XFILLER_0_187_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13733_ game.writer.tracker.frame\[218\] net845 net837 game.writer.tracker.frame\[217\]
+ vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_201_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10945_ game.CPU.applesa.ab.absxs.body_y\[28\] net533 vssd1 vssd1 vccd1 vccd1 _04835_
+ sky130_fd_sc_hd__or2_1
XANTENNA__16845__X _02619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19825__CLK clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19240_ clknet_leaf_16_clk _00071_ _00878_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.counter1.count\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_16452_ net186 net117 _02410_ _02406_ net1706 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[52\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_195_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13664_ _07534_ _07537_ net205 vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10876_ game.CPU.applesa.ab.apple_possible\[5\] game.CPU.applesa.ab.apple_possible\[6\]
+ game.CPU.applesa.ab.apple_possible\[7\] net551 vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__or4_1
XFILLER_0_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15403_ _01430_ _08906_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__and2b_1
XFILLER_0_213_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_356_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12615_ _06313_ _06315_ _06322_ _06491_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__a31o_1
XANTENNA__17389__A net1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19171_ clknet_leaf_4_clk _01290_ _00833_ vssd1 vssd1 vccd1 vccd1 game.CPU.randy.f1.a1.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_344_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16383_ net1927 net720 _02360_ vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[33\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__13946__A2 _03418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13595_ _07467_ _07468_ net515 vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__mux2_1
XANTENNA__17137__A2 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_225_Right_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11957__A1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18122_ net577 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11957__B2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_314_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15334_ _00029_ _08875_ _08876_ _08873_ _08874_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_152_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12546_ _06416_ _06417_ _06419_ _06422_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__or4b_1
XANTENNA__19975__CLK clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14525__B _07399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_289_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16896__A1 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18053_ net655 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15265_ _08816_ _08819_ _08820_ vssd1 vssd1 vccd1 vccd1 _08821_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09619__B game.CPU.applesa.ab.check_walls.above.walls\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12326__A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12477_ game.CPU.applesa.ab.absxs.body_x\[31\] net528 vssd1 vssd1 vccd1 vccd1 _06354_
+ sky130_fd_sc_hd__xnor2_1
X_17004_ _02328_ _02440_ net86 net728 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__o31a_1
XANTENNA__11230__A game.CPU.applesa.ab.absxs.body_y\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _02179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09378__A2 game.CPU.applesa.ab.check_walls.above.walls\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14216_ game.CPU.applesa.ab.absxs.body_x\[94\] net877 net861 game.CPU.applesa.ab.absxs.body_y\[93\]
+ _08089_ vssd1 vssd1 vccd1 vccd1 _08090_ sky130_fd_sc_hd__a221o_1
X_11428_ game.CPU.applesa.ab.check_walls.above.walls\[29\] net317 vssd1 vssd1 vccd1
+ vccd1 _05317_ sky130_fd_sc_hd__nand2_1
X_15196_ game.CPU.applesa.normal1.number\[4\] game.CPU.applesa.normal1.counter_flip
+ vssd1 vssd1 vccd1 vccd1 _08766_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_285_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12045__B net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16648__A1 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_284_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19205__CLK clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_286_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11359_ _05239_ _05241_ _05243_ _05247_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14147_ _08008_ _08013_ _07895_ vssd1 vssd1 vccd1 vccd1 _08021_ sky130_fd_sc_hd__o21a_1
XFILLER_0_158_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_228_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18013__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09635__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_265_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11884__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18955_ net1199 _00088_ _00626_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_33_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14078_ net1173 net857 game.CPU.applesa.ab.YMAX\[2\] net852 vssd1 vssd1 vccd1 vccd1
+ _07952_ sky130_fd_sc_hd__o22a_1
XFILLER_0_308_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13331__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_292_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13029_ _06894_ _06896_ _06899_ _06902_ net287 net240 vssd1 vssd1 vccd1 vccd1 _06903_
+ sky130_fd_sc_hd__mux4_1
X_17906_ net668 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__inv_2
XFILLER_0_184_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15075__C net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18886_ clknet_leaf_6_clk game.CPU.randy.f1.c1.innerCount\[16\] _00581_ vssd1 vssd1
+ vccd1 vccd1 game.CPU.randy.f1.c1.count\[16\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_280_Left_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19355__CLK clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1060 net1062 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_163_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17073__A1 _02267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1071 game.CPU.applesa.x\[0\] vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_280_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17837_ net182 _03163_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__nor2_1
XANTENNA__09550__A2 game.CPU.applesa.ab.absxs.body_x\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_206_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1082 net1083 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_8
Xfanout1093 net1095 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_8
XANTENNA__16468__A net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_351_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16820__A1 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17768_ _03121_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__inv_2
XFILLER_0_233_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09838__B1 game.CPU.applesa.ab.absxs.body_y\[107\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_178_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16719_ net1934 _02572_ _02574_ net109 vssd1 vssd1 vccd1 vccd1 game.writer.tracker.next_frame\[155\]
+ sky130_fd_sc_hd__a22o_1
X_19507_ clknet_leaf_14_clk game.writer.tracker.next_frame\[102\] net1282 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[102\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15091__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_297_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17699_ game.CPU.walls.rand_wall.count\[2\] game.CPU.walls.rand_wall.count\[1\] game.CPU.walls.rand_wall.count\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__and3_1
XFILLER_0_159_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19438_ clknet_leaf_43_clk game.writer.tracker.next_frame\[33\] net1303 vssd1 vssd1
+ vccd1 vccd1 game.writer.tracker.frame\[33\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_239_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_308_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16474__Y _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11660__A3 _05206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_252_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11124__B net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_340_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19369_ clknet_leaf_71_clk _01375_ _00950_ vssd1 vssd1 vccd1 vccd1 game.CPU.apple_location2\[2\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__12935__S net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13493__S0 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09122_ net1172 vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10963__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ game.CPU.applesa.ab.absxs.body_y\[76\] vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__inv_2
XFILLER_0_303_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_288_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout212_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_303_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_288_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 game.CPU.applesa.ab.absxs.body_y\[2\] vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_331_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold521 game.writer.tracker.frame\[4\] vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 game.writer.tracker.frame\[429\] vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16639__A1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_349_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold543 game.writer.tracker.frame\[422\] vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12373__B2 game.CPU.applesa.ab.absxs.body_y\[112\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold554 game.writer.tracker.frame\[80\] vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 game.writer.tracker.frame\[412\] vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17300__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14451__A game.CPU.applesa.ab.absxs.body_y\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1121_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 game.writer.tracker.frame\[386\] vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_268_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold587 game.writer.tracker.frame\[37\] vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1219_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09545__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold598 game.CPU.randy.f1.c1.count\[9\] vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_263_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09955_ _04172_ _04185_ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__nor2_1
XANTENNA__14170__B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout581_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_283_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout679_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_256_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09886_ net924 _03787_ _03707_ _03608_ _03545_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__o2111a_1
XANTENNA__17064__A1 _02438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09832__X _04075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_271_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10687__A1 game.CPU.applesa.ab.absxs.body_y\[102\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10687__B2 game.CPU.applesa.ab.absxs.body_y\[98\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16378__A net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_252_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout846_A _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_X net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_327_Right_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_358_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_339_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_358_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_352_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10730_ game.CPU.applesa.ab.absxs.body_y\[29\] net330 _04714_ net2053 vssd1 vssd1
+ vccd1 vccd1 _01052_ sky130_fd_sc_hd__a22o_1
XANTENNA__18872__CLK clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_314_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19998__CLK clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_354_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16825__B net143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_250_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_216_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11034__B net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10661_ game.CPU.applesa.ab.absxs.body_x\[26\] _04695_ _04698_ game.CPU.applesa.ab.absxs.body_x\[22\]
+ vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__a22o_1
XANTENNA__19764__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13484__S0 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17119__A2 _02524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11939__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16544__C _02393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11939__B2 net572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12400_ game.CPU.applesa.ab.absxs.body_x\[92\] net381 vssd1 vssd1 vccd1 vccd1 _06277_
+ sky130_fd_sc_hd__xnor2_1
X_13380_ net276 _07246_ net238 vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__o21a_1
X_10592_ _04173_ _04593_ _04589_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12600__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19197__Q game.CPU.walls.rand_wall.good_spot vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_341_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_334_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12331_ net528 vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.twoapples.absxs.next_head\[3\]
+ sky130_fd_sc_hd__inv_6
XANTENNA__17937__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10611__B2 net1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_259_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12262_ net786 net421 vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__or2_1
X_15050_ net1215 net1241 net812 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_188_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14353__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13787__S1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_267_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12364__A1 game.CPU.applesa.ab.absxs.body_y\[45\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_259_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11213_ _05094_ _05095_ _05100_ _05101_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__a22o_1
X_14001_ _07872_ _07873_ _07874_ vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__nor3b_1
XANTENNA__14999__C game.CPU.applesa.ab.check_walls.above.walls\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12193_ game.CPU.applesa.ab.check_walls.above.walls\[29\] net549 vssd1 vssd1 vccd1
+ vccd1 _06079_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_247_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_247_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput41 net41 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XANTENNA__19378__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
X_11144_ game.CPU.applesa.ab.absxs.body_y\[98\] net403 vssd1 vssd1 vccd1 vccd1 _05034_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__14080__B game.CPU.applesa.ab.check_walls.above.walls\[93\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18740_ clknet_leaf_8_clk _01157_ _00477_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_x\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_275_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15952_ game.CPU.applesa.ab.check_walls.above.walls\[27\] net462 vssd1 vssd1 vccd1
+ vccd1 _01964_ sky130_fd_sc_hd__nor2_1
X_11075_ game.CPU.applesa.ab.absxs.body_x\[40\] net324 vssd1 vssd1 vccd1 vccd1 _04965_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__13864__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17055__A1 _02423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_262_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10026_ _04233_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__inv_2
X_14903_ _08678_ _08679_ vssd1 vssd1 vccd1 vccd1 _08680_ sky130_fd_sc_hd__and2b_1
XANTENNA__11209__B net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18671_ clknet_leaf_10_clk _01088_ _00408_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.body_y\[101\]
+ sky130_fd_sc_hd__dfrtp_4
X_15883_ _01891_ _01892_ _01893_ _01894_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__or4_1
XANTENNA__16288__A net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_215_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16802__A1 _02487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17622_ game.CPU.kyle.L1.cnt_20ms\[13\] _03028_ net577 vssd1 vssd1 vccd1 vccd1 _03030_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__15605__A2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_188_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14834_ game.CPU.randy.f1.c1.count\[3\] _08632_ vssd1 vssd1 vccd1 vccd1 _08635_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_199_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_230_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17553_ _03219_ _00039_ _02835_ _02978_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a31o_1
X_14765_ game.CPU.randy.counter1.count\[10\] game.CPU.randy.counter1.count\[9\] _08583_
+ _08585_ vssd1 vssd1 vccd1 vccd1 _08586_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_316_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ _05192_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__and2_1
X_16504_ _02229_ _02400_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__nor2_2
XANTENNA__11225__A game.CPU.applesa.ab.absxs.body_y\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_156_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13716_ net202 _07585_ _07589_ net284 vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__o211a_1
X_10928_ net1166 net1168 game.CPU.applesa.ab.apple_possible\[4\] _04256_ _04809_ vssd1
+ vssd1 vccd1 vccd1 game.CPU.applesa.ab.absxs.next_head\[4\] sky130_fd_sc_hd__a311o_1
X_17484_ _02901_ _02902_ _02907_ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__and3_1
XFILLER_0_224_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14696_ game.CPU.randy.counter1.count1\[15\] _08499_ _08527_ vssd1 vssd1 vccd1 vccd1
+ _08535_ sky130_fd_sc_hd__a21bo_1
X_19223_ clknet_leaf_69_clk _01317_ _00862_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.apple_location\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_344_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_329_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16435_ game.writer.tracker.frame\[48\] _02395_ _02397_ net136 vssd1 vssd1 vccd1
+ vccd1 game.writer.tracker.next_frame\[48\] sky130_fd_sc_hd__a22o_1
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13647_ net513 _07517_ _07518_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__and3_1
XANTENNA__12755__S net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10859_ _03498_ game.CPU.randy.counter1.count1\[15\] vssd1 vssd1 vccd1 vccd1 _04762_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__14041__A1 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14041__B2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18008__A net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_17_Left_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19154_ net1187 _00197_ _00825_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[199\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09599__A2 game.CPU.applesa.ab.absxs.body_x\[75\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16366_ net197 _02347_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__nor2_4
X_13578_ net212 _07451_ net283 vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_288_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18105_ net632 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15317_ game.CPU.applesa.twomode.counter _08859_ _08860_ _08861_ _08862_ vssd1 vssd1
+ vccd1 vccd1 _08863_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19085_ net1178 _00122_ _00756_ vssd1 vssd1 vccd1 vccd1 game.CPU.applesa.ab.check_walls.above.walls\[130\]
+ sky130_fd_sc_hd__dfrtp_4
X_12529_ game.CPU.applesa.ab.absxs.body_x\[97\] net376 net368 game.CPU.applesa.ab.absxs.body_y\[99\]
+ _06405_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__a221o_1
X_16297_ net235 _02296_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__nor2_2
XFILLER_0_124_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_313_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18036_ net605 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__inv_2
XFILLER_0_340_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15541__A1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15248_ _00293_ _08808_ vssd1 vssd1 vccd1 vccd1 _08809_ sky130_fd_sc_hd__and2_4
XANTENNA__14344__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16470__B _02341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_297_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15179_ game.CPU.bodymain1.main.score\[5\] game.CPU.bodymain1.main.score\[4\] _04176_
+ _04581_ _04577_ vssd1 vssd1 vccd1 vccd1 _08755_ sky130_fd_sc_hd__a41o_1
XFILLER_0_319_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15086__B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 net309 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_272_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout319 game.CPU.applesa.ab.absxs.next_head\[2\] vssd1 vssd1 vccd1 vccd1 net319
+ sky130_fd_sc_hd__buf_6
X_19987_ clknet_leaf_44_clk _01411_ net1304 vssd1 vssd1 vccd1 vccd1 game.writer.updater.commands.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_26_Left_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18745__CLK clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ net1112 game.CPU.applesa.ab.check_walls.above.walls\[64\] vssd1 vssd1 vccd1
+ vccd1 _03983_ sky130_fd_sc_hd__xor2_1
XFILLER_0_185_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18938_ net1176 _00077_ vssd1 vssd1 vccd1 vccd1 game.CPU.walls.abc.number_out\[0\]
+ sky130_fd_sc_hd__dfxtp_1
.ends

